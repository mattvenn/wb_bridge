magic
tech sky130A
magscale 1 2
timestamp 1640939653
<< locali >>
rect 10977 77095 11011 78625
rect 10977 70907 11011 73525
rect 765 59143 799 69241
rect 11069 68935 11103 72437
rect 857 65127 891 66453
rect 949 65059 983 66113
rect 11161 65535 11195 72505
rect 11253 65807 11287 76789
rect 11437 74537 11471 77333
rect 11437 74503 11563 74537
rect 10977 65501 11195 65535
rect 949 64447 983 65025
rect 857 64413 949 64447
rect 857 62883 891 64413
rect 857 60095 891 62849
rect 765 55267 799 56389
rect 949 55539 983 64005
rect 765 53567 799 55233
rect 857 55505 983 55539
rect 857 53431 891 55505
rect 213 41531 247 44285
rect 673 42891 707 47685
rect 765 43843 799 48161
rect 857 40035 891 45509
rect 949 41803 983 55369
rect 10977 46699 11011 65501
rect 11069 58599 11103 62645
rect 11253 60737 11287 65637
rect 11161 60703 11287 60737
rect 11069 53567 11103 56661
rect 10977 42619 11011 46529
rect 3065 42007 3099 42177
rect 949 41769 1075 41803
rect 765 29019 799 36805
rect 857 30311 891 34493
rect 949 32351 983 41565
rect 1041 41531 1075 41769
rect 11069 36839 11103 53397
rect 11161 37927 11195 60703
rect 11253 52071 11287 55573
rect 11345 53431 11379 65705
rect 11253 34459 11287 51901
rect 11345 42143 11379 46665
rect 11437 41417 11471 65909
rect 11529 65127 11563 74503
rect 11621 61115 11655 65773
rect 11529 55403 11563 59381
rect 11621 49895 11655 57409
rect 11713 49419 11747 56865
rect 11805 50235 11839 58497
rect 11897 51935 11931 59109
rect 11345 41383 11471 41417
rect 11345 38471 11379 41383
rect 949 23307 983 28917
rect 10977 23239 11011 30685
rect 11069 24395 11103 31297
rect 11161 29767 11195 32861
rect 11253 23851 11287 31773
rect 10977 14943 11011 17153
rect 11069 16235 11103 19329
rect 10977 10251 11011 14365
rect 11069 10183 11103 16065
rect 11161 15623 11195 20893
rect 11161 9163 11195 13889
rect 11253 9367 11287 14977
<< viali >>
rect 10977 78625 11011 78659
rect 1409 77537 1443 77571
rect 1685 77537 1719 77571
rect 2881 77469 2915 77503
rect 3985 77469 4019 77503
rect 4629 77469 4663 77503
rect 9413 77469 9447 77503
rect 10057 77469 10091 77503
rect 2697 77333 2731 77367
rect 3801 77333 3835 77367
rect 4445 77333 4479 77367
rect 9229 77333 9263 77367
rect 9965 77333 9999 77367
rect 4445 77129 4479 77163
rect 9229 77129 9263 77163
rect 1593 77061 1627 77095
rect 1685 77061 1719 77095
rect 10057 77061 10091 77095
rect 10977 77061 11011 77095
rect 11437 77333 11471 77367
rect 1409 76993 1443 77027
rect 1829 76993 1863 77027
rect 2697 76993 2731 77027
rect 3341 76993 3375 77027
rect 3985 76993 4019 77027
rect 4629 76993 4663 77027
rect 9413 76993 9447 77027
rect 1961 76857 1995 76891
rect 2513 76789 2547 76823
rect 3157 76789 3191 76823
rect 3801 76789 3835 76823
rect 9965 76789 9999 76823
rect 11253 76789 11287 76823
rect 2421 76517 2455 76551
rect 3801 76517 3835 76551
rect 1869 76381 1903 76415
rect 2053 76381 2087 76415
rect 2242 76381 2276 76415
rect 3157 76381 3191 76415
rect 3985 76381 4019 76415
rect 10149 76381 10183 76415
rect 2145 76313 2179 76347
rect 2973 76245 3007 76279
rect 9965 76245 9999 76279
rect 1593 76041 1627 76075
rect 3433 76041 3467 76075
rect 9965 76041 9999 76075
rect 2513 75973 2547 76007
rect 2605 75973 2639 76007
rect 1409 75905 1443 75939
rect 2329 75905 2363 75939
rect 2702 75905 2736 75939
rect 3617 75905 3651 75939
rect 10149 75905 10183 75939
rect 2881 75701 2915 75735
rect 2421 75429 2455 75463
rect 1869 75293 1903 75327
rect 2053 75293 2087 75327
rect 2242 75293 2276 75327
rect 3157 75293 3191 75327
rect 10149 75293 10183 75327
rect 2145 75225 2179 75259
rect 2973 75157 3007 75191
rect 9965 75157 9999 75191
rect 2697 74885 2731 74919
rect 1409 74817 1443 74851
rect 2461 74817 2495 74851
rect 2605 74817 2639 74851
rect 2881 74817 2915 74851
rect 1593 74613 1627 74647
rect 2329 74613 2363 74647
rect 1409 74205 1443 74239
rect 10149 74205 10183 74239
rect 1593 74069 1627 74103
rect 9965 74069 9999 74103
rect 1869 73797 1903 73831
rect 1680 73729 1714 73763
rect 1777 73729 1811 73763
rect 2053 73729 2087 73763
rect 2697 73729 2731 73763
rect 10149 73729 10183 73763
rect 1501 73525 1535 73559
rect 2513 73525 2547 73559
rect 9965 73525 9999 73559
rect 10977 73525 11011 73559
rect 1680 73117 1714 73151
rect 1777 73117 1811 73151
rect 2032 73117 2066 73151
rect 2513 73117 2547 73151
rect 1869 73049 1903 73083
rect 1493 72981 1527 73015
rect 2697 72981 2731 73015
rect 2605 72709 2639 72743
rect 1409 72641 1443 72675
rect 2461 72641 2495 72675
rect 2697 72641 2731 72675
rect 2881 72641 2915 72675
rect 10149 72641 10183 72675
rect 1593 72437 1627 72471
rect 2329 72437 2363 72471
rect 9965 72437 9999 72471
rect 9965 72233 9999 72267
rect 1409 72029 1443 72063
rect 2053 72029 2087 72063
rect 10149 72029 10183 72063
rect 1593 71893 1627 71927
rect 2237 71893 2271 71927
rect 9965 71689 9999 71723
rect 1409 71553 1443 71587
rect 2237 71553 2271 71587
rect 10149 71553 10183 71587
rect 1593 71349 1627 71383
rect 2053 71349 2087 71383
rect 2789 71077 2823 71111
rect 1409 70941 1443 70975
rect 2237 70941 2271 70975
rect 2421 70941 2455 70975
rect 2610 70941 2644 70975
rect 11161 72505 11195 72539
rect 2513 70873 2547 70907
rect 10977 70873 11011 70907
rect 11069 72437 11103 72471
rect 1593 70805 1627 70839
rect 2513 70601 2547 70635
rect 9965 70601 9999 70635
rect 1593 70533 1627 70567
rect 1685 70533 1719 70567
rect 1409 70465 1443 70499
rect 1782 70465 1816 70499
rect 2697 70465 2731 70499
rect 10149 70465 10183 70499
rect 1961 70329 1995 70363
rect 1961 69989 1995 70023
rect 1409 69853 1443 69887
rect 1593 69853 1627 69887
rect 1782 69853 1816 69887
rect 2697 69853 2731 69887
rect 10149 69853 10183 69887
rect 1685 69785 1719 69819
rect 2513 69717 2547 69751
rect 9965 69717 9999 69751
rect 1593 69445 1627 69479
rect 1409 69377 1443 69411
rect 1685 69377 1719 69411
rect 1782 69377 1816 69411
rect 2697 69377 2731 69411
rect 3341 69377 3375 69411
rect 765 69241 799 69275
rect 1961 69173 1995 69207
rect 2513 69173 2547 69207
rect 3157 69173 3191 69207
rect 9965 68969 9999 69003
rect 11069 68901 11103 68935
rect 1409 68765 1443 68799
rect 2508 68765 2542 68799
rect 2605 68765 2639 68799
rect 2881 68765 2915 68799
rect 10149 68765 10183 68799
rect 2697 68697 2731 68731
rect 1593 68629 1627 68663
rect 2321 68629 2355 68663
rect 9965 68425 9999 68459
rect 2881 68357 2915 68391
rect 2973 68357 3007 68391
rect 1685 68289 1719 68323
rect 2697 68289 2731 68323
rect 3070 68289 3104 68323
rect 10149 68289 10183 68323
rect 1409 68221 1443 68255
rect 3249 68085 3283 68119
rect 1685 67745 1719 67779
rect 1409 67677 1443 67711
rect 1685 67201 1719 67235
rect 10149 67201 10183 67235
rect 1409 67133 1443 67167
rect 9965 66997 9999 67031
rect 1409 66589 1443 66623
rect 1685 66589 1719 66623
rect 2973 66589 3007 66623
rect 10149 66589 10183 66623
rect 857 66453 891 66487
rect 2789 66453 2823 66487
rect 9965 66453 9999 66487
rect 1593 66181 1627 66215
rect 2697 66181 2731 66215
rect 2789 66181 2823 66215
rect 857 65093 891 65127
rect 949 66113 983 66147
rect 1409 66113 1443 66147
rect 1685 66113 1719 66147
rect 1829 66113 1863 66147
rect 2513 66113 2547 66147
rect 2933 66113 2967 66147
rect 10149 66113 10183 66147
rect 1961 65977 1995 66011
rect 9965 65977 9999 66011
rect 3065 65909 3099 65943
rect 2145 65637 2179 65671
rect 11253 65773 11287 65807
rect 11437 65909 11471 65943
rect 11345 65705 11379 65739
rect 1409 65501 1443 65535
rect 2277 65501 2311 65535
rect 2421 65501 2455 65535
rect 2559 65501 2593 65535
rect 2697 65501 2731 65535
rect 3801 65501 3835 65535
rect 11253 65637 11287 65671
rect 1593 65365 1627 65399
rect 3985 65365 4019 65399
rect 1961 65161 1995 65195
rect 1593 65093 1627 65127
rect 1685 65093 1719 65127
rect 949 65025 983 65059
rect 1409 65025 1443 65059
rect 1777 65025 1811 65059
rect 2973 65025 3007 65059
rect 3249 65025 3283 65059
rect 3709 65025 3743 65059
rect 10149 65025 10183 65059
rect 3893 64889 3927 64923
rect 9965 64821 9999 64855
rect 1961 64549 1995 64583
rect 949 64413 983 64447
rect 1409 64413 1443 64447
rect 1593 64413 1627 64447
rect 1829 64413 1863 64447
rect 2513 64413 2547 64447
rect 10149 64413 10183 64447
rect 1685 64345 1719 64379
rect 2697 64277 2731 64311
rect 9965 64277 9999 64311
rect 857 62849 891 62883
rect 857 60061 891 60095
rect 949 64005 983 64039
rect 765 59109 799 59143
rect 765 56389 799 56423
rect 1685 63937 1719 63971
rect 2421 63937 2455 63971
rect 1501 63733 1535 63767
rect 2237 63733 2271 63767
rect 2329 63461 2363 63495
rect 1685 63325 1719 63359
rect 2145 63325 2179 63359
rect 2881 63325 2915 63359
rect 10149 63325 10183 63359
rect 1501 63189 1535 63223
rect 3065 63189 3099 63223
rect 9965 63189 9999 63223
rect 1593 62917 1627 62951
rect 1685 62917 1719 62951
rect 1409 62849 1443 62883
rect 1829 62849 1863 62883
rect 2881 62849 2915 62883
rect 3157 62849 3191 62883
rect 10149 62849 10183 62883
rect 1961 62713 1995 62747
rect 9965 62645 9999 62679
rect 2697 62305 2731 62339
rect 1685 62237 1719 62271
rect 2973 62237 3007 62271
rect 10149 62237 10183 62271
rect 1501 62101 1535 62135
rect 9965 62101 9999 62135
rect 1685 61761 1719 61795
rect 2421 61761 2455 61795
rect 2237 61625 2271 61659
rect 1501 61557 1535 61591
rect 1685 61149 1719 61183
rect 2421 61149 2455 61183
rect 2605 61149 2639 61183
rect 2789 61149 2823 61183
rect 10149 61149 10183 61183
rect 2697 61081 2731 61115
rect 1501 61013 1535 61047
rect 2973 61013 3007 61047
rect 9965 61013 9999 61047
rect 1685 60741 1719 60775
rect 1547 60673 1581 60707
rect 1777 60673 1811 60707
rect 1921 60673 1955 60707
rect 2605 60673 2639 60707
rect 10149 60673 10183 60707
rect 2789 60537 2823 60571
rect 2053 60469 2087 60503
rect 9965 60469 9999 60503
rect 2605 60197 2639 60231
rect 2053 60061 2087 60095
rect 2473 60061 2507 60095
rect 2237 59993 2271 60027
rect 2329 59993 2363 60027
rect 2329 59653 2363 59687
rect 2421 59653 2455 59687
rect 1685 59585 1719 59619
rect 2145 59585 2179 59619
rect 2565 59585 2599 59619
rect 3249 59585 3283 59619
rect 10149 59585 10183 59619
rect 3433 59449 3467 59483
rect 1501 59381 1535 59415
rect 2697 59381 2731 59415
rect 9965 59381 9999 59415
rect 2605 59177 2639 59211
rect 1961 59109 1995 59143
rect 1409 58973 1443 59007
rect 1593 58973 1627 59007
rect 1829 58973 1863 59007
rect 2789 58973 2823 59007
rect 10149 58973 10183 59007
rect 1685 58905 1719 58939
rect 9965 58837 9999 58871
rect 1869 58565 1903 58599
rect 1725 58497 1759 58531
rect 1961 58497 1995 58531
rect 2145 58497 2179 58531
rect 2605 58497 2639 58531
rect 9873 58497 9907 58531
rect 10149 58429 10183 58463
rect 1593 58293 1627 58327
rect 2789 58293 2823 58327
rect 1501 57885 1535 57919
rect 1921 57885 1955 57919
rect 2070 57885 2104 57919
rect 2605 57885 2639 57919
rect 3893 57885 3927 57919
rect 3985 57885 4019 57919
rect 1685 57817 1719 57851
rect 1777 57817 1811 57851
rect 2789 57749 2823 57783
rect 2973 57545 3007 57579
rect 1685 57409 1719 57443
rect 2421 57409 2455 57443
rect 2881 57409 2915 57443
rect 3065 57409 3099 57443
rect 9873 57409 9907 57443
rect 10149 57341 10183 57375
rect 2237 57273 2271 57307
rect 1501 57205 1535 57239
rect 3065 57001 3099 57035
rect 9873 56865 9907 56899
rect 1685 56797 1719 56831
rect 2421 56797 2455 56831
rect 2881 56797 2915 56831
rect 3065 56797 3099 56831
rect 3801 56797 3835 56831
rect 3985 56797 4019 56831
rect 10149 56797 10183 56831
rect 1501 56661 1535 56695
rect 2237 56661 2271 56695
rect 3893 56661 3927 56695
rect 2605 56389 2639 56423
rect 1685 56321 1719 56355
rect 2881 56321 2915 56355
rect 3341 56321 3375 56355
rect 3525 56321 3559 56355
rect 1501 56117 1535 56151
rect 3525 56117 3559 56151
rect 2973 55913 3007 55947
rect 1685 55709 1719 55743
rect 2145 55709 2179 55743
rect 3065 55709 3099 55743
rect 10149 55709 10183 55743
rect 1501 55573 1535 55607
rect 2329 55573 2363 55607
rect 9965 55573 9999 55607
rect 765 55233 799 55267
rect 765 53533 799 53567
rect 857 53397 891 53431
rect 949 55369 983 55403
rect 765 48161 799 48195
rect 673 47685 707 47719
rect 213 44285 247 44319
rect 765 43809 799 43843
rect 857 45509 891 45543
rect 673 42857 707 42891
rect 213 41497 247 41531
rect 1593 55301 1627 55335
rect 1685 55301 1719 55335
rect 3341 55301 3375 55335
rect 1409 55233 1443 55267
rect 1777 55233 1811 55267
rect 2605 55233 2639 55267
rect 10149 55233 10183 55267
rect 1961 55029 1995 55063
rect 9965 55029 9999 55063
rect 1685 54621 1719 54655
rect 2145 54621 2179 54655
rect 1501 54485 1535 54519
rect 2329 54485 2363 54519
rect 1685 54145 1719 54179
rect 2789 54145 2823 54179
rect 2973 54145 3007 54179
rect 9873 54145 9907 54179
rect 10057 54009 10091 54043
rect 1501 53941 1535 53975
rect 2973 53941 3007 53975
rect 2697 53737 2731 53771
rect 1978 53601 2012 53635
rect 1409 53533 1443 53567
rect 1593 53533 1627 53567
rect 1829 53533 1863 53567
rect 2513 53533 2547 53567
rect 2697 53533 2731 53567
rect 9873 53533 9907 53567
rect 1685 53465 1719 53499
rect 10057 53397 10091 53431
rect 1685 53057 1719 53091
rect 2145 53057 2179 53091
rect 2881 53057 2915 53091
rect 9873 53057 9907 53091
rect 3065 52921 3099 52955
rect 1501 52853 1535 52887
rect 2329 52853 2363 52887
rect 10057 52853 10091 52887
rect 2237 52649 2271 52683
rect 1685 52445 1719 52479
rect 2237 52445 2271 52479
rect 2421 52445 2455 52479
rect 1501 52309 1535 52343
rect 2513 52105 2547 52139
rect 1593 52037 1627 52071
rect 1685 52037 1719 52071
rect 1409 51969 1443 52003
rect 1777 51969 1811 52003
rect 2421 51969 2455 52003
rect 2605 51969 2639 52003
rect 3065 51969 3099 52003
rect 3249 51969 3283 52003
rect 9873 51969 9907 52003
rect 3157 51901 3191 51935
rect 1961 51833 1995 51867
rect 10057 51765 10091 51799
rect 1685 51357 1719 51391
rect 2421 51357 2455 51391
rect 2881 51357 2915 51391
rect 9873 51357 9907 51391
rect 1501 51221 1535 51255
rect 2237 51221 2271 51255
rect 3065 51221 3099 51255
rect 10057 51221 10091 51255
rect 3157 51017 3191 51051
rect 1685 50881 1719 50915
rect 3065 50881 3099 50915
rect 3249 50881 3283 50915
rect 1501 50677 1535 50711
rect 2605 50473 2639 50507
rect 3065 50473 3099 50507
rect 3985 50473 4019 50507
rect 1593 50269 1627 50303
rect 1685 50269 1719 50303
rect 1961 50269 1995 50303
rect 2421 50269 2455 50303
rect 2605 50269 2639 50303
rect 3065 50269 3099 50303
rect 3249 50269 3283 50303
rect 3801 50269 3835 50303
rect 3985 50269 4019 50303
rect 9873 50269 9907 50303
rect 1777 50201 1811 50235
rect 1409 50133 1443 50167
rect 10057 50133 10091 50167
rect 1685 49861 1719 49895
rect 1593 49793 1627 49827
rect 1777 49793 1811 49827
rect 1961 49793 1995 49827
rect 2421 49793 2455 49827
rect 9873 49793 9907 49827
rect 1409 49589 1443 49623
rect 2605 49589 2639 49623
rect 10057 49589 10091 49623
rect 1409 49181 1443 49215
rect 1685 49181 1719 49215
rect 1777 49181 1811 49215
rect 2421 49181 2455 49215
rect 3801 49181 3835 49215
rect 9873 49181 9907 49215
rect 1593 49113 1627 49147
rect 4077 49113 4111 49147
rect 1961 49045 1995 49079
rect 2605 49045 2639 49079
rect 10057 49045 10091 49079
rect 2237 48841 2271 48875
rect 1685 48705 1719 48739
rect 2421 48705 2455 48739
rect 1501 48501 1535 48535
rect 1685 48093 1719 48127
rect 2605 48093 2639 48127
rect 2789 48093 2823 48127
rect 9873 48093 9907 48127
rect 1501 47957 1535 47991
rect 2697 47957 2731 47991
rect 10057 47957 10091 47991
rect 2973 47753 3007 47787
rect 1685 47617 1719 47651
rect 2421 47617 2455 47651
rect 2881 47617 2915 47651
rect 3065 47617 3099 47651
rect 3525 47617 3559 47651
rect 3709 47617 3743 47651
rect 9873 47617 9907 47651
rect 3617 47549 3651 47583
rect 2237 47481 2271 47515
rect 1501 47413 1535 47447
rect 10057 47413 10091 47447
rect 2421 47209 2455 47243
rect 3065 47209 3099 47243
rect 1685 47005 1719 47039
rect 2237 47005 2271 47039
rect 2421 47005 2455 47039
rect 2881 47005 2915 47039
rect 3065 47005 3099 47039
rect 1501 46869 1535 46903
rect 11069 62645 11103 62679
rect 11069 58565 11103 58599
rect 11069 56661 11103 56695
rect 11069 53533 11103 53567
rect 10977 46665 11011 46699
rect 11069 53397 11103 53431
rect 1685 46529 1719 46563
rect 2513 46529 2547 46563
rect 2697 46529 2731 46563
rect 9873 46529 9907 46563
rect 10977 46529 11011 46563
rect 2697 46393 2731 46427
rect 10057 46393 10091 46427
rect 1501 46325 1535 46359
rect 1685 45917 1719 45951
rect 9873 45917 9907 45951
rect 1501 45781 1535 45815
rect 10057 45781 10091 45815
rect 1685 45441 1719 45475
rect 2329 45441 2363 45475
rect 1501 45237 1535 45271
rect 2145 45237 2179 45271
rect 1961 44965 1995 44999
rect 1777 44829 1811 44863
rect 1961 44829 1995 44863
rect 2513 44829 2547 44863
rect 9873 44829 9907 44863
rect 2697 44693 2731 44727
rect 10057 44693 10091 44727
rect 1501 44489 1535 44523
rect 1685 44353 1719 44387
rect 2145 44353 2179 44387
rect 3157 44353 3191 44387
rect 3617 44353 3651 44387
rect 3801 44353 3835 44387
rect 9873 44353 9907 44387
rect 3709 44285 3743 44319
rect 2329 44149 2363 44183
rect 2973 44149 3007 44183
rect 10057 44149 10091 44183
rect 1501 43809 1535 43843
rect 1593 43741 1627 43775
rect 1777 43741 1811 43775
rect 2605 43741 2639 43775
rect 3065 43741 3099 43775
rect 3249 43741 3283 43775
rect 9873 43741 9907 43775
rect 2421 43605 2455 43639
rect 3157 43605 3191 43639
rect 10057 43605 10091 43639
rect 3341 43401 3375 43435
rect 4629 43401 4663 43435
rect 1685 43333 1719 43367
rect 3985 43333 4019 43367
rect 1869 43265 1903 43299
rect 1961 43265 1995 43299
rect 2513 43265 2547 43299
rect 3249 43265 3283 43299
rect 3433 43265 3467 43299
rect 3893 43265 3927 43299
rect 4077 43265 4111 43299
rect 4537 43265 4571 43299
rect 4721 43265 4755 43299
rect 2697 43061 2731 43095
rect 1593 42857 1627 42891
rect 1409 42653 1443 42687
rect 1593 42653 1627 42687
rect 2145 42653 2179 42687
rect 2421 42653 2455 42687
rect 2881 42653 2915 42687
rect 3801 42653 3835 42687
rect 3985 42653 4019 42687
rect 9873 42653 9907 42687
rect 3893 42585 3927 42619
rect 10977 42585 11011 42619
rect 2145 42517 2179 42551
rect 3065 42517 3099 42551
rect 10057 42517 10091 42551
rect 3249 42313 3283 42347
rect 1685 42177 1719 42211
rect 2421 42177 2455 42211
rect 3065 42177 3099 42211
rect 3157 42177 3191 42211
rect 3341 42177 3375 42211
rect 9873 42177 9907 42211
rect 1501 41973 1535 42007
rect 2237 41973 2271 42007
rect 3065 41973 3099 42007
rect 10057 41973 10091 42007
rect 2973 41769 3007 41803
rect 857 40001 891 40035
rect 949 41565 983 41599
rect 765 36805 799 36839
rect 857 34493 891 34527
rect 1961 41633 1995 41667
rect 2145 41565 2179 41599
rect 2329 41565 2363 41599
rect 2789 41565 2823 41599
rect 2973 41565 3007 41599
rect 1041 41497 1075 41531
rect 1685 41089 1719 41123
rect 2421 41089 2455 41123
rect 2881 41089 2915 41123
rect 9873 41089 9907 41123
rect 3065 40953 3099 40987
rect 10057 40953 10091 40987
rect 1501 40885 1535 40919
rect 2237 40885 2271 40919
rect 2145 40681 2179 40715
rect 1685 40477 1719 40511
rect 2145 40477 2179 40511
rect 2329 40477 2363 40511
rect 9873 40477 9907 40511
rect 1501 40341 1535 40375
rect 10057 40341 10091 40375
rect 2237 40069 2271 40103
rect 1685 40001 1719 40035
rect 2145 40001 2179 40035
rect 2329 40001 2363 40035
rect 2881 40001 2915 40035
rect 3065 40001 3099 40035
rect 9873 40001 9907 40035
rect 3065 39865 3099 39899
rect 1501 39797 1535 39831
rect 10057 39797 10091 39831
rect 1593 39457 1627 39491
rect 1685 39389 1719 39423
rect 1961 39389 1995 39423
rect 2421 39389 2455 39423
rect 2605 39253 2639 39287
rect 1961 39049 1995 39083
rect 4077 39049 4111 39083
rect 1869 38913 1903 38947
rect 2789 38913 2823 38947
rect 3249 38913 3283 38947
rect 3985 38913 4019 38947
rect 4169 38913 4203 38947
rect 9873 38913 9907 38947
rect 2605 38709 2639 38743
rect 3433 38709 3467 38743
rect 10057 38709 10091 38743
rect 3157 38505 3191 38539
rect 2145 38369 2179 38403
rect 3893 38369 3927 38403
rect 1685 38301 1719 38335
rect 2237 38301 2271 38335
rect 2421 38301 2455 38335
rect 2973 38301 3007 38335
rect 3157 38301 3191 38335
rect 3801 38301 3835 38335
rect 3985 38301 4019 38335
rect 9873 38301 9907 38335
rect 1501 38165 1535 38199
rect 10057 38165 10091 38199
rect 2237 37961 2271 37995
rect 3249 37961 3283 37995
rect 1685 37825 1719 37859
rect 2237 37825 2271 37859
rect 2513 37825 2547 37859
rect 3065 37825 3099 37859
rect 3341 37825 3375 37859
rect 1501 37621 1535 37655
rect 2605 37281 2639 37315
rect 1501 37213 1535 37247
rect 1685 37213 1719 37247
rect 2513 37213 2547 37247
rect 2697 37213 2731 37247
rect 9873 37213 9907 37247
rect 1869 37145 1903 37179
rect 10057 37077 10091 37111
rect 11253 55573 11287 55607
rect 11345 53397 11379 53431
rect 11253 52037 11287 52071
rect 11161 37893 11195 37927
rect 11253 51901 11287 51935
rect 11069 36805 11103 36839
rect 1685 36737 1719 36771
rect 2145 36737 2179 36771
rect 2881 36737 2915 36771
rect 9873 36737 9907 36771
rect 3065 36601 3099 36635
rect 1501 36533 1535 36567
rect 2329 36533 2363 36567
rect 10057 36533 10091 36567
rect 3249 36329 3283 36363
rect 1869 36261 1903 36295
rect 1961 36125 1995 36159
rect 2145 36125 2179 36159
rect 3065 36125 3099 36159
rect 3249 36125 3283 36159
rect 9873 36125 9907 36159
rect 10057 35989 10091 36023
rect 2329 35785 2363 35819
rect 2145 35649 2179 35683
rect 2329 35649 2363 35683
rect 2881 35649 2915 35683
rect 3065 35513 3099 35547
rect 3985 35241 4019 35275
rect 2789 35173 2823 35207
rect 1961 35037 1995 35071
rect 2145 35037 2179 35071
rect 2789 35037 2823 35071
rect 3065 35037 3099 35071
rect 3801 35037 3835 35071
rect 3985 35037 4019 35071
rect 9873 35037 9907 35071
rect 2237 34969 2271 35003
rect 10057 34901 10091 34935
rect 3249 34697 3283 34731
rect 1869 34629 1903 34663
rect 1593 34561 1627 34595
rect 1685 34561 1719 34595
rect 2605 34561 2639 34595
rect 3065 34561 3099 34595
rect 9873 34561 9907 34595
rect 11345 46665 11379 46699
rect 11345 42109 11379 42143
rect 11529 65093 11563 65127
rect 11621 65773 11655 65807
rect 11621 61081 11655 61115
rect 11529 59381 11563 59415
rect 11897 59109 11931 59143
rect 11805 58497 11839 58531
rect 11529 55369 11563 55403
rect 11621 57409 11655 57443
rect 11621 49861 11655 49895
rect 11713 56865 11747 56899
rect 11897 51901 11931 51935
rect 11805 50201 11839 50235
rect 11713 49385 11747 49419
rect 11345 38437 11379 38471
rect 11253 34425 11287 34459
rect 2421 34357 2455 34391
rect 10057 34357 10091 34391
rect 1501 34153 1535 34187
rect 3065 34153 3099 34187
rect 1685 33949 1719 33983
rect 2145 33949 2179 33983
rect 2881 33949 2915 33983
rect 3065 33949 3099 33983
rect 2329 33813 2363 33847
rect 2973 33609 3007 33643
rect 1409 33473 1443 33507
rect 2145 33473 2179 33507
rect 2881 33473 2915 33507
rect 9873 33473 9907 33507
rect 10057 33337 10091 33371
rect 1593 33269 1627 33303
rect 2329 33269 2363 33303
rect 3985 33065 4019 33099
rect 3065 32997 3099 33031
rect 1409 32861 1443 32895
rect 2145 32861 2179 32895
rect 2881 32861 2915 32895
rect 3065 32861 3099 32895
rect 3801 32861 3835 32895
rect 3985 32861 4019 32895
rect 9873 32861 9907 32895
rect 11161 32861 11195 32895
rect 1593 32725 1627 32759
rect 2329 32725 2363 32759
rect 10057 32725 10091 32759
rect 2881 32521 2915 32555
rect 1685 32385 1719 32419
rect 2789 32385 2823 32419
rect 2973 32385 3007 32419
rect 949 32317 983 32351
rect 1501 32181 1535 32215
rect 2053 31977 2087 32011
rect 2697 31909 2731 31943
rect 10057 31909 10091 31943
rect 2053 31773 2087 31807
rect 2513 31773 2547 31807
rect 9873 31773 9907 31807
rect 2421 31433 2455 31467
rect 1593 31365 1627 31399
rect 1869 31297 1903 31331
rect 2605 31297 2639 31331
rect 9873 31297 9907 31331
rect 11069 31297 11103 31331
rect 10057 31093 10091 31127
rect 2053 30889 2087 30923
rect 2789 30889 2823 30923
rect 3801 30889 3835 30923
rect 2237 30685 2271 30719
rect 2881 30685 2915 30719
rect 3985 30685 4019 30719
rect 9413 30685 9447 30719
rect 9873 30685 9907 30719
rect 10977 30685 11011 30719
rect 10057 30549 10091 30583
rect 2421 30345 2455 30379
rect 3709 30345 3743 30379
rect 857 30277 891 30311
rect 1685 30209 1719 30243
rect 2237 30209 2271 30243
rect 2421 30209 2455 30243
rect 3065 30209 3099 30243
rect 3249 30209 3283 30243
rect 3893 30209 3927 30243
rect 1501 30073 1535 30107
rect 10149 30005 10183 30039
rect 1501 29801 1535 29835
rect 3801 29801 3835 29835
rect 3249 29733 3283 29767
rect 2237 29665 2271 29699
rect 1593 29597 1627 29631
rect 2329 29597 2363 29631
rect 2605 29597 2639 29631
rect 3065 29597 3099 29631
rect 3249 29597 3283 29631
rect 3985 29597 4019 29631
rect 1593 29257 1627 29291
rect 2513 29257 2547 29291
rect 3065 29257 3099 29291
rect 1409 29121 1443 29155
rect 2329 29121 2363 29155
rect 2513 29121 2547 29155
rect 3249 29121 3283 29155
rect 765 28985 799 29019
rect 949 28917 983 28951
rect 2329 28713 2363 28747
rect 3065 28713 3099 28747
rect 1777 28645 1811 28679
rect 1777 28509 1811 28543
rect 2421 28509 2455 28543
rect 2881 28509 2915 28543
rect 10149 28373 10183 28407
rect 1593 28169 1627 28203
rect 2237 28169 2271 28203
rect 1777 28033 1811 28067
rect 2421 28033 2455 28067
rect 2053 27557 2087 27591
rect 2789 27557 2823 27591
rect 4905 27489 4939 27523
rect 1409 27421 1443 27455
rect 2053 27421 2087 27455
rect 2973 27421 3007 27455
rect 4169 27421 4203 27455
rect 1593 27285 1627 27319
rect 10149 27285 10183 27319
rect 2973 27081 3007 27115
rect 1593 27013 1627 27047
rect 1869 26945 1903 26979
rect 2513 26945 2547 26979
rect 3157 26945 3191 26979
rect 2421 26809 2455 26843
rect 1501 26537 1535 26571
rect 2881 26537 2915 26571
rect 2145 26469 2179 26503
rect 10149 26401 10183 26435
rect 1685 26333 1719 26367
rect 2237 26333 2271 26367
rect 3065 26333 3099 26367
rect 2237 25993 2271 26027
rect 2697 25993 2731 26027
rect 1409 25857 1443 25891
rect 2053 25857 2087 25891
rect 2881 25857 2915 25891
rect 1593 25653 1627 25687
rect 1961 25449 1995 25483
rect 10149 25449 10183 25483
rect 1961 25245 1995 25279
rect 2605 25245 2639 25279
rect 2421 25109 2455 25143
rect 1409 24769 1443 24803
rect 2145 24769 2179 24803
rect 2973 24769 3007 24803
rect 10149 24769 10183 24803
rect 2237 24701 2271 24735
rect 2789 24633 2823 24667
rect 1593 24565 1627 24599
rect 1685 24361 1719 24395
rect 2881 24361 2915 24395
rect 1869 24157 1903 24191
rect 2697 24157 2731 24191
rect 2881 24157 2915 24191
rect 3985 24157 4019 24191
rect 3801 24021 3835 24055
rect 3801 23817 3835 23851
rect 1409 23681 1443 23715
rect 2053 23681 2087 23715
rect 2329 23681 2363 23715
rect 2973 23681 3007 23715
rect 3249 23681 3283 23715
rect 3709 23681 3743 23715
rect 3893 23681 3927 23715
rect 9873 23681 9907 23715
rect 2421 23613 2455 23647
rect 2973 23545 3007 23579
rect 1593 23477 1627 23511
rect 10057 23477 10091 23511
rect 949 23273 983 23307
rect 9505 23273 9539 23307
rect 10149 23273 10183 23307
rect 11161 29733 11195 29767
rect 11253 31773 11287 31807
rect 11069 24361 11103 24395
rect 11253 23817 11287 23851
rect 1961 23205 1995 23239
rect 3985 23205 4019 23239
rect 10977 23205 11011 23239
rect 1685 23069 1719 23103
rect 1961 23069 1995 23103
rect 2789 23069 2823 23103
rect 3801 23069 3835 23103
rect 3985 23069 4019 23103
rect 9321 23069 9355 23103
rect 3065 23001 3099 23035
rect 1501 22729 1535 22763
rect 3893 22729 3927 22763
rect 1409 22593 1443 22627
rect 2421 22593 2455 22627
rect 4077 22593 4111 22627
rect 9873 22593 9907 22627
rect 2789 22525 2823 22559
rect 10057 22457 10091 22491
rect 2973 22185 3007 22219
rect 1593 22049 1627 22083
rect 1685 21981 1719 22015
rect 2329 21981 2363 22015
rect 2421 21981 2455 22015
rect 3157 21981 3191 22015
rect 9229 21981 9263 22015
rect 9873 21981 9907 22015
rect 2421 21845 2455 21879
rect 9413 21845 9447 21879
rect 10057 21845 10091 21879
rect 2973 21641 3007 21675
rect 1409 21505 1443 21539
rect 2513 21505 2547 21539
rect 9873 21505 9907 21539
rect 1593 21301 1627 21335
rect 2605 21301 2639 21335
rect 10057 21301 10091 21335
rect 2237 21097 2271 21131
rect 3065 21097 3099 21131
rect 9873 21097 9907 21131
rect 3801 21029 3835 21063
rect 1685 20893 1719 20927
rect 2421 20893 2455 20927
rect 2881 20893 2915 20927
rect 3985 20893 4019 20927
rect 10057 20893 10091 20927
rect 11161 20893 11195 20927
rect 1593 20757 1627 20791
rect 3157 20553 3191 20587
rect 2053 20417 2087 20451
rect 2697 20417 2731 20451
rect 3341 20417 3375 20451
rect 9873 20417 9907 20451
rect 2513 20281 2547 20315
rect 10057 20281 10091 20315
rect 1961 20213 1995 20247
rect 1869 20009 1903 20043
rect 1869 19805 1903 19839
rect 2513 19805 2547 19839
rect 3157 19805 3191 19839
rect 9873 19805 9907 19839
rect 2329 19669 2363 19703
rect 2973 19669 3007 19703
rect 10057 19669 10091 19703
rect 9873 19465 9907 19499
rect 1869 19329 1903 19363
rect 2329 19329 2363 19363
rect 10057 19329 10091 19363
rect 11069 19329 11103 19363
rect 1869 19193 1903 19227
rect 2513 19125 2547 19159
rect 1777 18921 1811 18955
rect 9413 18921 9447 18955
rect 3065 18785 3099 18819
rect 1777 18717 1811 18751
rect 2421 18717 2455 18751
rect 3985 18717 4019 18751
rect 9229 18717 9263 18751
rect 9873 18717 9907 18751
rect 3801 18581 3835 18615
rect 10057 18581 10091 18615
rect 1685 18377 1719 18411
rect 2421 18377 2455 18411
rect 9413 18377 9447 18411
rect 2605 18309 2639 18343
rect 2789 18309 2823 18343
rect 1777 18241 1811 18275
rect 3433 18241 3467 18275
rect 9229 18241 9263 18275
rect 9873 18241 9907 18275
rect 3249 18037 3283 18071
rect 10057 18037 10091 18071
rect 1961 17833 1995 17867
rect 3801 17833 3835 17867
rect 2605 17765 2639 17799
rect 2053 17629 2087 17663
rect 2513 17629 2547 17663
rect 3985 17629 4019 17663
rect 9873 17629 9907 17663
rect 10057 17493 10091 17527
rect 9965 17289 9999 17323
rect 1409 17153 1443 17187
rect 2237 17153 2271 17187
rect 2881 17153 2915 17187
rect 10149 17153 10183 17187
rect 10977 17153 11011 17187
rect 1593 16949 1627 16983
rect 2053 16949 2087 16983
rect 2697 16949 2731 16983
rect 2145 16541 2179 16575
rect 2789 16541 2823 16575
rect 9229 16541 9263 16575
rect 9873 16541 9907 16575
rect 2053 16473 2087 16507
rect 2605 16405 2639 16439
rect 9413 16405 9447 16439
rect 10057 16405 10091 16439
rect 1961 16201 1995 16235
rect 2605 16201 2639 16235
rect 1501 16065 1535 16099
rect 1777 16065 1811 16099
rect 2421 16065 2455 16099
rect 2513 16065 2547 16099
rect 9873 16065 9907 16099
rect 1685 15997 1719 16031
rect 2789 15997 2823 16031
rect 1777 15861 1811 15895
rect 2513 15861 2547 15895
rect 10057 15861 10091 15895
rect 1501 15657 1535 15691
rect 9965 15657 9999 15691
rect 2697 15589 2731 15623
rect 1409 15453 1443 15487
rect 1593 15453 1627 15487
rect 2237 15453 2271 15487
rect 2881 15453 2915 15487
rect 10149 15453 10183 15487
rect 2053 15317 2087 15351
rect 1869 15113 1903 15147
rect 2973 15113 3007 15147
rect 1777 15045 1811 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2513 14977 2547 15011
rect 2789 14977 2823 15011
rect 9873 14977 9907 15011
rect 11069 16201 11103 16235
rect 2605 14909 2639 14943
rect 10977 14909 11011 14943
rect 11069 16065 11103 16099
rect 10057 14841 10091 14875
rect 1961 14773 1995 14807
rect 2513 14773 2547 14807
rect 1409 14569 1443 14603
rect 1869 14569 1903 14603
rect 2329 14569 2363 14603
rect 1777 14433 1811 14467
rect 1593 14365 1627 14399
rect 2513 14365 2547 14399
rect 3157 14365 3191 14399
rect 3985 14365 4019 14399
rect 9873 14365 9907 14399
rect 10977 14365 11011 14399
rect 1869 14297 1903 14331
rect 2973 14229 3007 14263
rect 3801 14229 3835 14263
rect 10057 14229 10091 14263
rect 1961 14025 1995 14059
rect 2881 14025 2915 14059
rect 9413 14025 9447 14059
rect 1869 13889 1903 13923
rect 2697 13889 2731 13923
rect 2881 13889 2915 13923
rect 9229 13889 9263 13923
rect 9873 13889 9907 13923
rect 10057 13685 10091 13719
rect 2973 13413 3007 13447
rect 1685 13345 1719 13379
rect 1409 13277 1443 13311
rect 2789 13209 2823 13243
rect 2789 12937 2823 12971
rect 1685 12801 1719 12835
rect 2973 12801 3007 12835
rect 9873 12801 9907 12835
rect 1409 12733 1443 12767
rect 10057 12597 10091 12631
rect 2789 12393 2823 12427
rect 1685 12257 1719 12291
rect 1409 12189 1443 12223
rect 2973 12189 3007 12223
rect 3801 12189 3835 12223
rect 9873 12189 9907 12223
rect 3985 12053 4019 12087
rect 10057 12053 10091 12087
rect 2789 11849 2823 11883
rect 1685 11713 1719 11747
rect 2973 11713 3007 11747
rect 3433 11713 3467 11747
rect 4077 11713 4111 11747
rect 1409 11645 1443 11679
rect 3617 11509 3651 11543
rect 4261 11509 4295 11543
rect 3985 11237 4019 11271
rect 10057 11237 10091 11271
rect 1685 11169 1719 11203
rect 1409 11101 1443 11135
rect 2697 11101 2731 11135
rect 3801 11101 3835 11135
rect 9873 11101 9907 11135
rect 2881 10965 2915 10999
rect 3433 10693 3467 10727
rect 1685 10625 1719 10659
rect 2973 10625 3007 10659
rect 3249 10625 3283 10659
rect 9873 10625 9907 10659
rect 1409 10557 1443 10591
rect 10057 10421 10091 10455
rect 9965 10217 9999 10251
rect 10977 10217 11011 10251
rect 11161 15589 11195 15623
rect 11253 14977 11287 15011
rect 9505 10149 9539 10183
rect 11069 10149 11103 10183
rect 11161 13889 11195 13923
rect 1685 10081 1719 10115
rect 1409 10013 1443 10047
rect 2697 10013 2731 10047
rect 9321 10013 9355 10047
rect 10149 10013 10183 10047
rect 2881 9877 2915 9911
rect 2789 9673 2823 9707
rect 2900 9605 2934 9639
rect 1685 9537 1719 9571
rect 2697 9537 2731 9571
rect 3065 9537 3099 9571
rect 9229 9537 9263 9571
rect 9873 9537 9907 9571
rect 1409 9469 1443 9503
rect 2789 9401 2823 9435
rect 10057 9401 10091 9435
rect 9413 9333 9447 9367
rect 11253 9333 11287 9367
rect 2421 9129 2455 9163
rect 3249 9129 3283 9163
rect 9413 9129 9447 9163
rect 11161 9129 11195 9163
rect 1869 8925 1903 8959
rect 2605 8925 2639 8959
rect 3065 8925 3099 8959
rect 9229 8925 9263 8959
rect 9873 8925 9907 8959
rect 1685 8789 1719 8823
rect 10057 8789 10091 8823
rect 1593 8585 1627 8619
rect 2329 8585 2363 8619
rect 3709 8585 3743 8619
rect 1409 8449 1443 8483
rect 2145 8449 2179 8483
rect 2881 8449 2915 8483
rect 3525 8449 3559 8483
rect 9873 8449 9907 8483
rect 3065 8313 3099 8347
rect 10057 8245 10091 8279
rect 3985 8041 4019 8075
rect 1685 7905 1719 7939
rect 1409 7837 1443 7871
rect 2697 7837 2731 7871
rect 3801 7837 3835 7871
rect 2881 7701 2915 7735
rect 2789 7497 2823 7531
rect 1869 7429 1903 7463
rect 1961 7361 1995 7395
rect 2605 7361 2639 7395
rect 3341 7361 3375 7395
rect 3525 7361 3559 7395
rect 9873 7361 9907 7395
rect 3525 7157 3559 7191
rect 10057 7157 10091 7191
rect 1409 6749 1443 6783
rect 2605 6749 2639 6783
rect 9873 6749 9907 6783
rect 1593 6613 1627 6647
rect 2789 6613 2823 6647
rect 10057 6613 10091 6647
rect 1593 6409 1627 6443
rect 2237 6409 2271 6443
rect 3525 6409 3559 6443
rect 1409 6273 1443 6307
rect 2053 6273 2087 6307
rect 2697 6273 2731 6307
rect 3341 6273 3375 6307
rect 2881 6137 2915 6171
rect 1593 5865 1627 5899
rect 1409 5661 1443 5695
rect 2329 5661 2363 5695
rect 9873 5661 9907 5695
rect 2513 5525 2547 5559
rect 10057 5525 10091 5559
rect 1593 5321 1627 5355
rect 2237 5253 2271 5287
rect 1409 5185 1443 5219
rect 2329 5185 2363 5219
rect 2789 5185 2823 5219
rect 2973 5185 3007 5219
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4077 5185 4111 5219
rect 4261 5185 4295 5219
rect 9873 5185 9907 5219
rect 2973 4981 3007 5015
rect 3617 4981 3651 5015
rect 4261 4981 4295 5015
rect 10057 4981 10091 5015
rect 2237 4777 2271 4811
rect 3801 4777 3835 4811
rect 2789 4709 2823 4743
rect 2237 4573 2271 4607
rect 2881 4573 2915 4607
rect 3985 4573 4019 4607
rect 9873 4573 9907 4607
rect 10057 4437 10091 4471
rect 2053 4165 2087 4199
rect 1593 4097 1627 4131
rect 2329 4097 2363 4131
rect 2513 4097 2547 4131
rect 3249 4097 3283 4131
rect 3433 4097 3467 4131
rect 3893 4097 3927 4131
rect 4077 4097 4111 4131
rect 1501 4029 1535 4063
rect 3433 3961 3467 3995
rect 4077 3893 4111 3927
rect 3801 3689 3835 3723
rect 2145 3485 2179 3519
rect 2697 3485 2731 3519
rect 3985 3485 4019 3519
rect 9873 3485 9907 3519
rect 2605 3349 2639 3383
rect 10057 3349 10091 3383
rect 2237 3145 2271 3179
rect 3433 3145 3467 3179
rect 4077 3145 4111 3179
rect 1685 3009 1719 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3617 3009 3651 3043
rect 4261 3009 4295 3043
rect 9137 3009 9171 3043
rect 9873 3009 9907 3043
rect 2973 2873 3007 2907
rect 1501 2805 1535 2839
rect 9321 2805 9355 2839
rect 10057 2805 10091 2839
rect 1593 2601 1627 2635
rect 2697 2601 2731 2635
rect 3801 2601 3835 2635
rect 4445 2601 4479 2635
rect 5089 2601 5123 2635
rect 2237 2533 2271 2567
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 5273 2397 5307 2431
rect 9137 2397 9171 2431
rect 9873 2397 9907 2431
rect 9321 2261 9355 2295
rect 10057 2261 10091 2295
<< metal1 >>
rect 10962 78656 10968 78668
rect 10923 78628 10968 78656
rect 10962 78616 10968 78628
rect 11020 78616 11026 78668
rect 2774 78072 2780 78124
rect 2832 78112 2838 78124
rect 4614 78112 4620 78124
rect 2832 78084 4620 78112
rect 2832 78072 2838 78084
rect 4614 78072 4620 78084
rect 4672 78072 4678 78124
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5845 77818
rect 5897 77766 5909 77818
rect 5961 77766 5973 77818
rect 6025 77766 6037 77818
rect 6089 77766 6101 77818
rect 6153 77766 9109 77818
rect 9161 77766 9173 77818
rect 9225 77766 9237 77818
rect 9289 77766 9301 77818
rect 9353 77766 9365 77818
rect 9417 77766 10856 77818
rect 1104 77744 10856 77766
rect 1394 77568 1400 77580
rect 1355 77540 1400 77568
rect 1394 77528 1400 77540
rect 1452 77528 1458 77580
rect 1673 77571 1731 77577
rect 1673 77537 1685 77571
rect 1719 77568 1731 77571
rect 3602 77568 3608 77580
rect 1719 77540 3608 77568
rect 1719 77537 1731 77540
rect 1673 77531 1731 77537
rect 3602 77528 3608 77540
rect 3660 77528 3666 77580
rect 2869 77503 2927 77509
rect 2869 77469 2881 77503
rect 2915 77500 2927 77503
rect 2958 77500 2964 77512
rect 2915 77472 2964 77500
rect 2915 77469 2927 77472
rect 2869 77463 2927 77469
rect 2958 77460 2964 77472
rect 3016 77460 3022 77512
rect 3970 77500 3976 77512
rect 3931 77472 3976 77500
rect 3970 77460 3976 77472
rect 4028 77460 4034 77512
rect 4062 77460 4068 77512
rect 4120 77500 4126 77512
rect 4617 77503 4675 77509
rect 4617 77500 4629 77503
rect 4120 77472 4629 77500
rect 4120 77460 4126 77472
rect 4617 77469 4629 77472
rect 4663 77469 4675 77503
rect 9398 77500 9404 77512
rect 9359 77472 9404 77500
rect 4617 77463 4675 77469
rect 9398 77460 9404 77472
rect 9456 77460 9462 77512
rect 10042 77500 10048 77512
rect 10003 77472 10048 77500
rect 10042 77460 10048 77472
rect 10100 77460 10106 77512
rect 2130 77324 2136 77376
rect 2188 77364 2194 77376
rect 2685 77367 2743 77373
rect 2685 77364 2697 77367
rect 2188 77336 2697 77364
rect 2188 77324 2194 77336
rect 2685 77333 2697 77336
rect 2731 77333 2743 77367
rect 3786 77364 3792 77376
rect 3747 77336 3792 77364
rect 2685 77327 2743 77333
rect 3786 77324 3792 77336
rect 3844 77324 3850 77376
rect 3878 77324 3884 77376
rect 3936 77364 3942 77376
rect 4433 77367 4491 77373
rect 4433 77364 4445 77367
rect 3936 77336 4445 77364
rect 3936 77324 3942 77336
rect 4433 77333 4445 77336
rect 4479 77333 4491 77367
rect 4433 77327 4491 77333
rect 5258 77324 5264 77376
rect 5316 77364 5322 77376
rect 9217 77367 9275 77373
rect 9217 77364 9229 77367
rect 5316 77336 9229 77364
rect 5316 77324 5322 77336
rect 9217 77333 9229 77336
rect 9263 77333 9275 77367
rect 9217 77327 9275 77333
rect 9953 77367 10011 77373
rect 9953 77333 9965 77367
rect 9999 77364 10011 77367
rect 11425 77367 11483 77373
rect 11425 77364 11437 77367
rect 9999 77336 11437 77364
rect 9999 77333 10011 77336
rect 9953 77327 10011 77333
rect 11425 77333 11437 77336
rect 11471 77333 11483 77367
rect 11425 77327 11483 77333
rect 1104 77274 10856 77296
rect 1104 77222 4213 77274
rect 4265 77222 4277 77274
rect 4329 77222 4341 77274
rect 4393 77222 4405 77274
rect 4457 77222 4469 77274
rect 4521 77222 7477 77274
rect 7529 77222 7541 77274
rect 7593 77222 7605 77274
rect 7657 77222 7669 77274
rect 7721 77222 7733 77274
rect 7785 77222 10856 77274
rect 1104 77200 10856 77222
rect 4433 77163 4491 77169
rect 4433 77160 4445 77163
rect 1596 77132 4445 77160
rect 1596 77101 1624 77132
rect 4433 77129 4445 77132
rect 4479 77129 4491 77163
rect 9217 77163 9275 77169
rect 9217 77160 9229 77163
rect 4433 77123 4491 77129
rect 6886 77132 9229 77160
rect 1581 77095 1639 77101
rect 1581 77061 1593 77095
rect 1627 77061 1639 77095
rect 1581 77055 1639 77061
rect 1673 77095 1731 77101
rect 1673 77061 1685 77095
rect 1719 77092 1731 77095
rect 6886 77092 6914 77132
rect 9217 77129 9229 77132
rect 9263 77129 9275 77163
rect 9217 77123 9275 77129
rect 1719 77064 6914 77092
rect 10045 77095 10103 77101
rect 1719 77061 1731 77064
rect 1673 77055 1731 77061
rect 10045 77061 10057 77095
rect 10091 77092 10103 77095
rect 10965 77095 11023 77101
rect 10965 77092 10977 77095
rect 10091 77064 10977 77092
rect 10091 77061 10103 77064
rect 10045 77055 10103 77061
rect 10965 77061 10977 77064
rect 11011 77061 11023 77095
rect 10965 77055 11023 77061
rect 1394 77024 1400 77036
rect 1355 76996 1400 77024
rect 1394 76984 1400 76996
rect 1452 76984 1458 77036
rect 1817 77027 1875 77033
rect 1817 76993 1829 77027
rect 1863 77024 1875 77027
rect 2222 77024 2228 77036
rect 1863 76996 2228 77024
rect 1863 76993 1875 76996
rect 1817 76987 1875 76993
rect 2222 76984 2228 76996
rect 2280 76984 2286 77036
rect 2685 77027 2743 77033
rect 2685 76993 2697 77027
rect 2731 77024 2743 77027
rect 2958 77024 2964 77036
rect 2731 76996 2964 77024
rect 2731 76993 2743 76996
rect 2685 76987 2743 76993
rect 2958 76984 2964 76996
rect 3016 76984 3022 77036
rect 3326 77024 3332 77036
rect 3287 76996 3332 77024
rect 3326 76984 3332 76996
rect 3384 76984 3390 77036
rect 3418 76984 3424 77036
rect 3476 77024 3482 77036
rect 3973 77027 4031 77033
rect 3973 77024 3985 77027
rect 3476 76996 3985 77024
rect 3476 76984 3482 76996
rect 3973 76993 3985 76996
rect 4019 76993 4031 77027
rect 4614 77024 4620 77036
rect 4575 76996 4620 77024
rect 3973 76987 4031 76993
rect 4614 76984 4620 76996
rect 4672 76984 4678 77036
rect 9401 77027 9459 77033
rect 9401 76993 9413 77027
rect 9447 77024 9459 77027
rect 9490 77024 9496 77036
rect 9447 76996 9496 77024
rect 9447 76993 9459 76996
rect 9401 76987 9459 76993
rect 9490 76984 9496 76996
rect 9548 76984 9554 77036
rect 1949 76891 2007 76897
rect 1949 76857 1961 76891
rect 1995 76888 2007 76891
rect 5534 76888 5540 76900
rect 1995 76860 5540 76888
rect 1995 76857 2007 76860
rect 1949 76851 2007 76857
rect 5534 76848 5540 76860
rect 5592 76848 5598 76900
rect 2406 76780 2412 76832
rect 2464 76820 2470 76832
rect 2501 76823 2559 76829
rect 2501 76820 2513 76823
rect 2464 76792 2513 76820
rect 2464 76780 2470 76792
rect 2501 76789 2513 76792
rect 2547 76789 2559 76823
rect 2501 76783 2559 76789
rect 3050 76780 3056 76832
rect 3108 76820 3114 76832
rect 3145 76823 3203 76829
rect 3145 76820 3157 76823
rect 3108 76792 3157 76820
rect 3108 76780 3114 76792
rect 3145 76789 3157 76792
rect 3191 76789 3203 76823
rect 3145 76783 3203 76789
rect 3234 76780 3240 76832
rect 3292 76820 3298 76832
rect 3789 76823 3847 76829
rect 3789 76820 3801 76823
rect 3292 76792 3801 76820
rect 3292 76780 3298 76792
rect 3789 76789 3801 76792
rect 3835 76789 3847 76823
rect 3789 76783 3847 76789
rect 9953 76823 10011 76829
rect 9953 76789 9965 76823
rect 9999 76820 10011 76823
rect 11241 76823 11299 76829
rect 11241 76820 11253 76823
rect 9999 76792 11253 76820
rect 9999 76789 10011 76792
rect 9953 76783 10011 76789
rect 11241 76789 11253 76792
rect 11287 76789 11299 76823
rect 11241 76783 11299 76789
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5845 76730
rect 5897 76678 5909 76730
rect 5961 76678 5973 76730
rect 6025 76678 6037 76730
rect 6089 76678 6101 76730
rect 6153 76678 9109 76730
rect 9161 76678 9173 76730
rect 9225 76678 9237 76730
rect 9289 76678 9301 76730
rect 9353 76678 9365 76730
rect 9417 76678 10856 76730
rect 1104 76656 10856 76678
rect 106 76508 112 76560
rect 164 76548 170 76560
rect 2409 76551 2467 76557
rect 2409 76548 2421 76551
rect 164 76520 2421 76548
rect 164 76508 170 76520
rect 2409 76517 2421 76520
rect 2455 76517 2467 76551
rect 2409 76511 2467 76517
rect 3789 76551 3847 76557
rect 3789 76517 3801 76551
rect 3835 76517 3847 76551
rect 3789 76511 3847 76517
rect 3804 76480 3832 76511
rect 2056 76452 3832 76480
rect 1394 76372 1400 76424
rect 1452 76412 1458 76424
rect 1857 76415 1915 76421
rect 1857 76412 1869 76415
rect 1452 76384 1869 76412
rect 1452 76372 1458 76384
rect 1857 76381 1869 76384
rect 1903 76412 1915 76415
rect 1946 76412 1952 76424
rect 1903 76384 1952 76412
rect 1903 76381 1915 76384
rect 1857 76375 1915 76381
rect 1946 76372 1952 76384
rect 2004 76372 2010 76424
rect 2056 76421 2084 76452
rect 2041 76415 2099 76421
rect 2041 76381 2053 76415
rect 2087 76381 2099 76415
rect 2041 76375 2099 76381
rect 2222 76372 2228 76424
rect 2280 76421 2286 76424
rect 2280 76412 2288 76421
rect 3142 76412 3148 76424
rect 2280 76384 2325 76412
rect 3103 76384 3148 76412
rect 2280 76375 2288 76384
rect 2280 76372 2286 76375
rect 3142 76372 3148 76384
rect 3200 76372 3206 76424
rect 3510 76372 3516 76424
rect 3568 76412 3574 76424
rect 3973 76415 4031 76421
rect 3973 76412 3985 76415
rect 3568 76384 3985 76412
rect 3568 76372 3574 76384
rect 3973 76381 3985 76384
rect 4019 76381 4031 76415
rect 10134 76412 10140 76424
rect 10095 76384 10140 76412
rect 3973 76375 4031 76381
rect 10134 76372 10140 76384
rect 10192 76372 10198 76424
rect 2133 76347 2191 76353
rect 2133 76313 2145 76347
rect 2179 76344 2191 76347
rect 5258 76344 5264 76356
rect 2179 76316 5264 76344
rect 2179 76313 2191 76316
rect 2133 76307 2191 76313
rect 5258 76304 5264 76316
rect 5316 76304 5322 76356
rect 2961 76279 3019 76285
rect 2961 76245 2973 76279
rect 3007 76276 3019 76279
rect 3418 76276 3424 76288
rect 3007 76248 3424 76276
rect 3007 76245 3019 76248
rect 2961 76239 3019 76245
rect 3418 76236 3424 76248
rect 3476 76236 3482 76288
rect 9950 76276 9956 76288
rect 9911 76248 9956 76276
rect 9950 76236 9956 76248
rect 10008 76236 10014 76288
rect 1104 76186 10856 76208
rect 1104 76134 4213 76186
rect 4265 76134 4277 76186
rect 4329 76134 4341 76186
rect 4393 76134 4405 76186
rect 4457 76134 4469 76186
rect 4521 76134 7477 76186
rect 7529 76134 7541 76186
rect 7593 76134 7605 76186
rect 7657 76134 7669 76186
rect 7721 76134 7733 76186
rect 7785 76134 10856 76186
rect 1104 76112 10856 76134
rect 1581 76075 1639 76081
rect 1581 76041 1593 76075
rect 1627 76072 1639 76075
rect 1762 76072 1768 76084
rect 1627 76044 1768 76072
rect 1627 76041 1639 76044
rect 1581 76035 1639 76041
rect 1762 76032 1768 76044
rect 1820 76032 1826 76084
rect 3234 76072 3240 76084
rect 2516 76044 3240 76072
rect 2516 76013 2544 76044
rect 3234 76032 3240 76044
rect 3292 76032 3298 76084
rect 3326 76032 3332 76084
rect 3384 76072 3390 76084
rect 3421 76075 3479 76081
rect 3421 76072 3433 76075
rect 3384 76044 3433 76072
rect 3384 76032 3390 76044
rect 3421 76041 3433 76044
rect 3467 76041 3479 76075
rect 9953 76075 10011 76081
rect 9953 76072 9965 76075
rect 3421 76035 3479 76041
rect 6886 76044 9965 76072
rect 2501 76007 2559 76013
rect 2501 75973 2513 76007
rect 2547 75973 2559 76007
rect 2501 75967 2559 75973
rect 2593 76007 2651 76013
rect 2593 75973 2605 76007
rect 2639 76004 2651 76007
rect 6886 76004 6914 76044
rect 9953 76041 9965 76044
rect 9999 76041 10011 76075
rect 9953 76035 10011 76041
rect 2639 75976 6914 76004
rect 2639 75973 2651 75976
rect 2593 75967 2651 75973
rect 1397 75939 1455 75945
rect 1397 75905 1409 75939
rect 1443 75936 1455 75939
rect 1486 75936 1492 75948
rect 1443 75908 1492 75936
rect 1443 75905 1455 75908
rect 1397 75899 1455 75905
rect 1486 75896 1492 75908
rect 1544 75896 1550 75948
rect 1946 75896 1952 75948
rect 2004 75936 2010 75948
rect 2317 75939 2375 75945
rect 2317 75936 2329 75939
rect 2004 75908 2329 75936
rect 2004 75896 2010 75908
rect 2317 75905 2329 75908
rect 2363 75905 2375 75939
rect 2317 75899 2375 75905
rect 2690 75939 2748 75945
rect 2690 75905 2702 75939
rect 2736 75905 2748 75939
rect 2690 75899 2748 75905
rect 2222 75828 2228 75880
rect 2280 75868 2286 75880
rect 2705 75868 2733 75899
rect 3602 75896 3608 75948
rect 3660 75936 3666 75948
rect 10137 75939 10195 75945
rect 3660 75908 3705 75936
rect 3660 75896 3666 75908
rect 10137 75905 10149 75939
rect 10183 75936 10195 75939
rect 10183 75908 10272 75936
rect 10183 75905 10195 75908
rect 10137 75899 10195 75905
rect 10244 75880 10272 75908
rect 2280 75840 2733 75868
rect 2280 75828 2286 75840
rect 10226 75828 10232 75880
rect 10284 75828 10290 75880
rect 3234 75760 3240 75812
rect 3292 75800 3298 75812
rect 3510 75800 3516 75812
rect 3292 75772 3516 75800
rect 3292 75760 3298 75772
rect 3510 75760 3516 75772
rect 3568 75760 3574 75812
rect 2869 75735 2927 75741
rect 2869 75701 2881 75735
rect 2915 75732 2927 75735
rect 3970 75732 3976 75744
rect 2915 75704 3976 75732
rect 2915 75701 2927 75704
rect 2869 75695 2927 75701
rect 3970 75692 3976 75704
rect 4028 75692 4034 75744
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5845 75642
rect 5897 75590 5909 75642
rect 5961 75590 5973 75642
rect 6025 75590 6037 75642
rect 6089 75590 6101 75642
rect 6153 75590 9109 75642
rect 9161 75590 9173 75642
rect 9225 75590 9237 75642
rect 9289 75590 9301 75642
rect 9353 75590 9365 75642
rect 9417 75590 10856 75642
rect 1104 75568 10856 75590
rect 2409 75463 2467 75469
rect 2409 75429 2421 75463
rect 2455 75460 2467 75463
rect 8294 75460 8300 75472
rect 2455 75432 8300 75460
rect 2455 75429 2467 75432
rect 2409 75423 2467 75429
rect 8294 75420 8300 75432
rect 8352 75420 8358 75472
rect 3878 75392 3884 75404
rect 2056 75364 3884 75392
rect 1857 75327 1915 75333
rect 1857 75293 1869 75327
rect 1903 75324 1915 75327
rect 1946 75324 1952 75336
rect 1903 75296 1952 75324
rect 1903 75293 1915 75296
rect 1857 75287 1915 75293
rect 1946 75284 1952 75296
rect 2004 75284 2010 75336
rect 2056 75333 2084 75364
rect 3878 75352 3884 75364
rect 3936 75352 3942 75404
rect 2041 75327 2099 75333
rect 2041 75293 2053 75327
rect 2087 75293 2099 75327
rect 2041 75287 2099 75293
rect 2222 75284 2228 75336
rect 2280 75333 2286 75336
rect 2280 75324 2288 75333
rect 3142 75324 3148 75336
rect 2280 75296 2325 75324
rect 3103 75296 3148 75324
rect 2280 75287 2288 75296
rect 2280 75284 2286 75287
rect 3142 75284 3148 75296
rect 3200 75284 3206 75336
rect 9950 75324 9956 75336
rect 6886 75296 9956 75324
rect 2133 75259 2191 75265
rect 2133 75225 2145 75259
rect 2179 75256 2191 75259
rect 6886 75256 6914 75296
rect 9950 75284 9956 75296
rect 10008 75284 10014 75336
rect 10134 75324 10140 75336
rect 10095 75296 10140 75324
rect 10134 75284 10140 75296
rect 10192 75284 10198 75336
rect 2179 75228 6914 75256
rect 2179 75225 2191 75228
rect 2133 75219 2191 75225
rect 2958 75188 2964 75200
rect 2919 75160 2964 75188
rect 2958 75148 2964 75160
rect 3016 75148 3022 75200
rect 9950 75188 9956 75200
rect 9911 75160 9956 75188
rect 9950 75148 9956 75160
rect 10008 75148 10014 75200
rect 1104 75098 10856 75120
rect 1104 75046 4213 75098
rect 4265 75046 4277 75098
rect 4329 75046 4341 75098
rect 4393 75046 4405 75098
rect 4457 75046 4469 75098
rect 4521 75046 7477 75098
rect 7529 75046 7541 75098
rect 7593 75046 7605 75098
rect 7657 75046 7669 75098
rect 7721 75046 7733 75098
rect 7785 75046 10856 75098
rect 1104 75024 10856 75046
rect 2685 74919 2743 74925
rect 2685 74885 2697 74919
rect 2731 74916 2743 74919
rect 3786 74916 3792 74928
rect 2731 74888 3792 74916
rect 2731 74885 2743 74888
rect 2685 74879 2743 74885
rect 3786 74876 3792 74888
rect 3844 74876 3850 74928
rect 1394 74848 1400 74860
rect 1355 74820 1400 74848
rect 1394 74808 1400 74820
rect 1452 74808 1458 74860
rect 1670 74808 1676 74860
rect 1728 74848 1734 74860
rect 2222 74848 2228 74860
rect 1728 74820 2228 74848
rect 1728 74808 1734 74820
rect 2222 74808 2228 74820
rect 2280 74848 2286 74860
rect 2449 74851 2507 74857
rect 2449 74848 2461 74851
rect 2280 74820 2461 74848
rect 2280 74808 2286 74820
rect 2449 74817 2461 74820
rect 2495 74817 2507 74851
rect 2449 74811 2507 74817
rect 2593 74851 2651 74857
rect 2593 74817 2605 74851
rect 2639 74817 2651 74851
rect 2593 74811 2651 74817
rect 2869 74851 2927 74857
rect 2869 74817 2881 74851
rect 2915 74848 2927 74851
rect 3142 74848 3148 74860
rect 2915 74820 3148 74848
rect 2915 74817 2927 74820
rect 2869 74811 2927 74817
rect 2608 74780 2636 74811
rect 3142 74808 3148 74820
rect 3200 74808 3206 74860
rect 9950 74780 9956 74792
rect 2608 74752 9956 74780
rect 9950 74740 9956 74752
rect 10008 74740 10014 74792
rect 1578 74644 1584 74656
rect 1539 74616 1584 74644
rect 1578 74604 1584 74616
rect 1636 74604 1642 74656
rect 2317 74647 2375 74653
rect 2317 74613 2329 74647
rect 2363 74644 2375 74647
rect 5626 74644 5632 74656
rect 2363 74616 5632 74644
rect 2363 74613 2375 74616
rect 2317 74607 2375 74613
rect 5626 74604 5632 74616
rect 5684 74604 5690 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5845 74554
rect 5897 74502 5909 74554
rect 5961 74502 5973 74554
rect 6025 74502 6037 74554
rect 6089 74502 6101 74554
rect 6153 74502 9109 74554
rect 9161 74502 9173 74554
rect 9225 74502 9237 74554
rect 9289 74502 9301 74554
rect 9353 74502 9365 74554
rect 9417 74502 10856 74554
rect 1104 74480 10856 74502
rect 1394 74236 1400 74248
rect 1355 74208 1400 74236
rect 1394 74196 1400 74208
rect 1452 74196 1458 74248
rect 10134 74236 10140 74248
rect 10095 74208 10140 74236
rect 10134 74196 10140 74208
rect 10192 74196 10198 74248
rect 1486 74060 1492 74112
rect 1544 74100 1550 74112
rect 1581 74103 1639 74109
rect 1581 74100 1593 74103
rect 1544 74072 1593 74100
rect 1544 74060 1550 74072
rect 1581 74069 1593 74072
rect 1627 74069 1639 74103
rect 9950 74100 9956 74112
rect 9911 74072 9956 74100
rect 1581 74063 1639 74069
rect 9950 74060 9956 74072
rect 10008 74060 10014 74112
rect 1104 74010 10856 74032
rect 1104 73958 4213 74010
rect 4265 73958 4277 74010
rect 4329 73958 4341 74010
rect 4393 73958 4405 74010
rect 4457 73958 4469 74010
rect 4521 73958 7477 74010
rect 7529 73958 7541 74010
rect 7593 73958 7605 74010
rect 7657 73958 7669 74010
rect 7721 73958 7733 74010
rect 7785 73958 10856 74010
rect 1104 73936 10856 73958
rect 1857 73831 1915 73837
rect 1857 73797 1869 73831
rect 1903 73828 1915 73831
rect 2958 73828 2964 73840
rect 1903 73800 2964 73828
rect 1903 73797 1915 73800
rect 1857 73791 1915 73797
rect 2958 73788 2964 73800
rect 3016 73788 3022 73840
rect 1670 73769 1676 73772
rect 1668 73760 1676 73769
rect 1631 73732 1676 73760
rect 1668 73723 1676 73732
rect 1670 73720 1676 73723
rect 1728 73720 1734 73772
rect 1765 73763 1823 73769
rect 1765 73729 1777 73763
rect 1811 73729 1823 73763
rect 1765 73723 1823 73729
rect 1780 73692 1808 73723
rect 1946 73720 1952 73772
rect 2004 73760 2010 73772
rect 2041 73763 2099 73769
rect 2041 73760 2053 73763
rect 2004 73732 2053 73760
rect 2004 73720 2010 73732
rect 2041 73729 2053 73732
rect 2087 73760 2099 73763
rect 2222 73760 2228 73772
rect 2087 73732 2228 73760
rect 2087 73729 2099 73732
rect 2041 73723 2099 73729
rect 2222 73720 2228 73732
rect 2280 73720 2286 73772
rect 2685 73763 2743 73769
rect 2685 73729 2697 73763
rect 2731 73760 2743 73763
rect 2774 73760 2780 73772
rect 2731 73732 2780 73760
rect 2731 73729 2743 73732
rect 2685 73723 2743 73729
rect 2774 73720 2780 73732
rect 2832 73720 2838 73772
rect 10134 73760 10140 73772
rect 10095 73732 10140 73760
rect 10134 73720 10140 73732
rect 10192 73720 10198 73772
rect 9858 73692 9864 73704
rect 1780 73664 9864 73692
rect 9858 73652 9864 73664
rect 9916 73652 9922 73704
rect 566 73516 572 73568
rect 624 73556 630 73568
rect 1489 73559 1547 73565
rect 1489 73556 1501 73559
rect 624 73528 1501 73556
rect 624 73516 630 73528
rect 1489 73525 1501 73528
rect 1535 73525 1547 73559
rect 1489 73519 1547 73525
rect 1946 73516 1952 73568
rect 2004 73556 2010 73568
rect 2501 73559 2559 73565
rect 2501 73556 2513 73559
rect 2004 73528 2513 73556
rect 2004 73516 2010 73528
rect 2501 73525 2513 73528
rect 2547 73525 2559 73559
rect 2501 73519 2559 73525
rect 9953 73559 10011 73565
rect 9953 73525 9965 73559
rect 9999 73556 10011 73559
rect 10965 73559 11023 73565
rect 10965 73556 10977 73559
rect 9999 73528 10977 73556
rect 9999 73525 10011 73528
rect 9953 73519 10011 73525
rect 10965 73525 10977 73528
rect 11011 73525 11023 73559
rect 10965 73519 11023 73525
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5845 73466
rect 5897 73414 5909 73466
rect 5961 73414 5973 73466
rect 6025 73414 6037 73466
rect 6089 73414 6101 73466
rect 6153 73414 9109 73466
rect 9161 73414 9173 73466
rect 9225 73414 9237 73466
rect 9289 73414 9301 73466
rect 9353 73414 9365 73466
rect 9417 73414 10856 73466
rect 1104 73392 10856 73414
rect 2222 73216 2228 73228
rect 2135 73188 2228 73216
rect 1670 73157 1676 73160
rect 1668 73148 1676 73157
rect 1631 73120 1676 73148
rect 1668 73111 1676 73120
rect 1670 73108 1676 73111
rect 1728 73108 1734 73160
rect 1765 73151 1823 73157
rect 1765 73117 1777 73151
rect 1811 73148 1823 73151
rect 2020 73151 2078 73157
rect 1811 73120 1992 73148
rect 1811 73117 1823 73120
rect 1765 73111 1823 73117
rect 1854 73080 1860 73092
rect 1815 73052 1860 73080
rect 1854 73040 1860 73052
rect 1912 73040 1918 73092
rect 1964 73080 1992 73120
rect 2020 73117 2032 73151
rect 2066 73144 2078 73151
rect 2148 73144 2176 73188
rect 2222 73176 2228 73188
rect 2280 73216 2286 73228
rect 2958 73216 2964 73228
rect 2280 73188 2964 73216
rect 2280 73176 2286 73188
rect 2958 73176 2964 73188
rect 3016 73216 3022 73228
rect 3142 73216 3148 73228
rect 3016 73188 3148 73216
rect 3016 73176 3022 73188
rect 3142 73176 3148 73188
rect 3200 73176 3206 73228
rect 2066 73117 2176 73144
rect 2020 73116 2176 73117
rect 2501 73151 2559 73157
rect 2501 73117 2513 73151
rect 2547 73148 2559 73151
rect 2774 73148 2780 73160
rect 2547 73120 2780 73148
rect 2547 73117 2559 73120
rect 2020 73111 2078 73116
rect 2501 73111 2559 73117
rect 2774 73108 2780 73120
rect 2832 73108 2838 73160
rect 4062 73080 4068 73092
rect 1964 73052 4068 73080
rect 4062 73040 4068 73052
rect 4120 73040 4126 73092
rect 1481 73015 1539 73021
rect 1481 72981 1493 73015
rect 1527 73012 1539 73015
rect 2222 73012 2228 73024
rect 1527 72984 2228 73012
rect 1527 72981 1539 72984
rect 1481 72975 1539 72981
rect 2222 72972 2228 72984
rect 2280 72972 2286 73024
rect 2498 72972 2504 73024
rect 2556 73012 2562 73024
rect 2685 73015 2743 73021
rect 2685 73012 2697 73015
rect 2556 72984 2697 73012
rect 2556 72972 2562 72984
rect 2685 72981 2697 72984
rect 2731 72981 2743 73015
rect 2685 72975 2743 72981
rect 1104 72922 10856 72944
rect 1104 72870 4213 72922
rect 4265 72870 4277 72922
rect 4329 72870 4341 72922
rect 4393 72870 4405 72922
rect 4457 72870 4469 72922
rect 4521 72870 7477 72922
rect 7529 72870 7541 72922
rect 7593 72870 7605 72922
rect 7657 72870 7669 72922
rect 7721 72870 7733 72922
rect 7785 72870 10856 72922
rect 1104 72848 10856 72870
rect 1854 72768 1860 72820
rect 1912 72808 1918 72820
rect 3326 72808 3332 72820
rect 1912 72780 3332 72808
rect 1912 72768 1918 72780
rect 3326 72768 3332 72780
rect 3384 72768 3390 72820
rect 2593 72743 2651 72749
rect 2593 72709 2605 72743
rect 2639 72740 2651 72743
rect 9950 72740 9956 72752
rect 2639 72712 9956 72740
rect 2639 72709 2651 72712
rect 2593 72703 2651 72709
rect 9950 72700 9956 72712
rect 10008 72700 10014 72752
rect 1394 72672 1400 72684
rect 1355 72644 1400 72672
rect 1394 72632 1400 72644
rect 1452 72632 1458 72684
rect 1670 72632 1676 72684
rect 1728 72672 1734 72684
rect 2314 72672 2320 72684
rect 1728 72644 2320 72672
rect 1728 72632 1734 72644
rect 2314 72632 2320 72644
rect 2372 72672 2378 72684
rect 2449 72675 2507 72681
rect 2449 72672 2461 72675
rect 2372 72644 2461 72672
rect 2372 72632 2378 72644
rect 2449 72641 2461 72644
rect 2495 72641 2507 72675
rect 2449 72635 2507 72641
rect 2685 72675 2743 72681
rect 2685 72641 2697 72675
rect 2731 72641 2743 72675
rect 2685 72635 2743 72641
rect 2869 72675 2927 72681
rect 2869 72641 2881 72675
rect 2915 72672 2927 72675
rect 2958 72672 2964 72684
rect 2915 72644 2964 72672
rect 2915 72641 2927 72644
rect 2869 72635 2927 72641
rect 2700 72604 2728 72635
rect 2958 72632 2964 72644
rect 3016 72632 3022 72684
rect 10134 72672 10140 72684
rect 10095 72644 10140 72672
rect 10134 72632 10140 72644
rect 10192 72632 10198 72684
rect 3050 72604 3056 72616
rect 2700 72576 3056 72604
rect 3050 72564 3056 72576
rect 3108 72564 3114 72616
rect 4062 72564 4068 72616
rect 4120 72604 4126 72616
rect 9950 72604 9956 72616
rect 4120 72576 9956 72604
rect 4120 72564 4126 72576
rect 9950 72564 9956 72576
rect 10008 72564 10014 72616
rect 2222 72496 2228 72548
rect 2280 72536 2286 72548
rect 8386 72536 8392 72548
rect 2280 72508 8392 72536
rect 2280 72496 2286 72508
rect 8386 72496 8392 72508
rect 8444 72496 8450 72548
rect 11149 72539 11207 72545
rect 11149 72536 11161 72539
rect 8956 72508 11161 72536
rect 1581 72471 1639 72477
rect 1581 72437 1593 72471
rect 1627 72468 1639 72471
rect 1670 72468 1676 72480
rect 1627 72440 1676 72468
rect 1627 72437 1639 72440
rect 1581 72431 1639 72437
rect 1670 72428 1676 72440
rect 1728 72428 1734 72480
rect 2317 72471 2375 72477
rect 2317 72437 2329 72471
rect 2363 72468 2375 72471
rect 8956 72468 8984 72508
rect 11149 72505 11161 72508
rect 11195 72505 11207 72539
rect 11149 72499 11207 72505
rect 2363 72440 8984 72468
rect 9953 72471 10011 72477
rect 2363 72437 2375 72440
rect 2317 72431 2375 72437
rect 9953 72437 9965 72471
rect 9999 72468 10011 72471
rect 11057 72471 11115 72477
rect 11057 72468 11069 72471
rect 9999 72440 11069 72468
rect 9999 72437 10011 72440
rect 9953 72431 10011 72437
rect 11057 72437 11069 72440
rect 11103 72437 11115 72471
rect 11057 72431 11115 72437
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5845 72378
rect 5897 72326 5909 72378
rect 5961 72326 5973 72378
rect 6025 72326 6037 72378
rect 6089 72326 6101 72378
rect 6153 72326 9109 72378
rect 9161 72326 9173 72378
rect 9225 72326 9237 72378
rect 9289 72326 9301 72378
rect 9353 72326 9365 72378
rect 9417 72326 10856 72378
rect 1104 72304 10856 72326
rect 9950 72264 9956 72276
rect 9911 72236 9956 72264
rect 9950 72224 9956 72236
rect 10008 72224 10014 72276
rect 1210 72020 1216 72072
rect 1268 72060 1274 72072
rect 1397 72063 1455 72069
rect 1397 72060 1409 72063
rect 1268 72032 1409 72060
rect 1268 72020 1274 72032
rect 1397 72029 1409 72032
rect 1443 72029 1455 72063
rect 2038 72060 2044 72072
rect 1999 72032 2044 72060
rect 1397 72023 1455 72029
rect 2038 72020 2044 72032
rect 2096 72020 2102 72072
rect 10134 72060 10140 72072
rect 10095 72032 10140 72060
rect 10134 72020 10140 72032
rect 10192 72020 10198 72072
rect 1486 71884 1492 71936
rect 1544 71924 1550 71936
rect 1581 71927 1639 71933
rect 1581 71924 1593 71927
rect 1544 71896 1593 71924
rect 1544 71884 1550 71896
rect 1581 71893 1593 71896
rect 1627 71893 1639 71927
rect 1581 71887 1639 71893
rect 2225 71927 2283 71933
rect 2225 71893 2237 71927
rect 2271 71924 2283 71927
rect 2314 71924 2320 71936
rect 2271 71896 2320 71924
rect 2271 71893 2283 71896
rect 2225 71887 2283 71893
rect 2314 71884 2320 71896
rect 2372 71884 2378 71936
rect 1104 71834 10856 71856
rect 1104 71782 4213 71834
rect 4265 71782 4277 71834
rect 4329 71782 4341 71834
rect 4393 71782 4405 71834
rect 4457 71782 4469 71834
rect 4521 71782 7477 71834
rect 7529 71782 7541 71834
rect 7593 71782 7605 71834
rect 7657 71782 7669 71834
rect 7721 71782 7733 71834
rect 7785 71782 10856 71834
rect 1104 71760 10856 71782
rect 2038 71680 2044 71732
rect 2096 71720 2102 71732
rect 2222 71720 2228 71732
rect 2096 71692 2228 71720
rect 2096 71680 2102 71692
rect 2222 71680 2228 71692
rect 2280 71680 2286 71732
rect 9858 71680 9864 71732
rect 9916 71720 9922 71732
rect 9953 71723 10011 71729
rect 9953 71720 9965 71723
rect 9916 71692 9965 71720
rect 9916 71680 9922 71692
rect 9953 71689 9965 71692
rect 9999 71689 10011 71723
rect 9953 71683 10011 71689
rect 1302 71544 1308 71596
rect 1360 71584 1366 71596
rect 1397 71587 1455 71593
rect 1397 71584 1409 71587
rect 1360 71556 1409 71584
rect 1360 71544 1366 71556
rect 1397 71553 1409 71556
rect 1443 71553 1455 71587
rect 2222 71584 2228 71596
rect 2183 71556 2228 71584
rect 1397 71547 1455 71553
rect 2222 71544 2228 71556
rect 2280 71544 2286 71596
rect 10134 71584 10140 71596
rect 10095 71556 10140 71584
rect 10134 71544 10140 71556
rect 10192 71544 10198 71596
rect 1581 71383 1639 71389
rect 1581 71349 1593 71383
rect 1627 71380 1639 71383
rect 1854 71380 1860 71392
rect 1627 71352 1860 71380
rect 1627 71349 1639 71352
rect 1581 71343 1639 71349
rect 1854 71340 1860 71352
rect 1912 71340 1918 71392
rect 2041 71383 2099 71389
rect 2041 71349 2053 71383
rect 2087 71380 2099 71383
rect 2222 71380 2228 71392
rect 2087 71352 2228 71380
rect 2087 71349 2099 71352
rect 2041 71343 2099 71349
rect 2222 71340 2228 71352
rect 2280 71340 2286 71392
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5845 71290
rect 5897 71238 5909 71290
rect 5961 71238 5973 71290
rect 6025 71238 6037 71290
rect 6089 71238 6101 71290
rect 6153 71238 9109 71290
rect 9161 71238 9173 71290
rect 9225 71238 9237 71290
rect 9289 71238 9301 71290
rect 9353 71238 9365 71290
rect 9417 71238 10856 71290
rect 1104 71216 10856 71238
rect 2777 71111 2835 71117
rect 2777 71077 2789 71111
rect 2823 71108 2835 71111
rect 5074 71108 5080 71120
rect 2823 71080 5080 71108
rect 2823 71077 2835 71080
rect 2777 71071 2835 71077
rect 5074 71068 5080 71080
rect 5132 71068 5138 71120
rect 2038 71000 2044 71052
rect 2096 71040 2102 71052
rect 2096 71012 2636 71040
rect 2096 71000 2102 71012
rect 2608 70984 2636 71012
rect 1394 70972 1400 70984
rect 1355 70944 1400 70972
rect 1394 70932 1400 70944
rect 1452 70932 1458 70984
rect 2225 70975 2283 70981
rect 2225 70941 2237 70975
rect 2271 70941 2283 70975
rect 2406 70972 2412 70984
rect 2367 70944 2412 70972
rect 2225 70935 2283 70941
rect 1210 70864 1216 70916
rect 1268 70904 1274 70916
rect 2240 70904 2268 70935
rect 2406 70932 2412 70944
rect 2464 70932 2470 70984
rect 2590 70932 2596 70984
rect 2648 70981 2654 70984
rect 2648 70972 2656 70981
rect 2648 70944 2693 70972
rect 2648 70935 2656 70944
rect 2648 70932 2654 70935
rect 1268 70876 2268 70904
rect 1268 70864 1274 70876
rect 1581 70839 1639 70845
rect 1581 70805 1593 70839
rect 1627 70836 1639 70839
rect 2038 70836 2044 70848
rect 1627 70808 2044 70836
rect 1627 70805 1639 70808
rect 1581 70799 1639 70805
rect 2038 70796 2044 70808
rect 2096 70796 2102 70848
rect 2240 70836 2268 70876
rect 2501 70907 2559 70913
rect 2501 70873 2513 70907
rect 2547 70904 2559 70907
rect 10965 70907 11023 70913
rect 10965 70904 10977 70907
rect 2547 70876 10977 70904
rect 2547 70873 2559 70876
rect 2501 70867 2559 70873
rect 10965 70873 10977 70876
rect 11011 70873 11023 70907
rect 10965 70867 11023 70873
rect 2958 70836 2964 70848
rect 2240 70808 2964 70836
rect 2958 70796 2964 70808
rect 3016 70796 3022 70848
rect 1104 70746 10856 70768
rect 1104 70694 4213 70746
rect 4265 70694 4277 70746
rect 4329 70694 4341 70746
rect 4393 70694 4405 70746
rect 4457 70694 4469 70746
rect 4521 70694 7477 70746
rect 7529 70694 7541 70746
rect 7593 70694 7605 70746
rect 7657 70694 7669 70746
rect 7721 70694 7733 70746
rect 7785 70694 10856 70746
rect 1104 70672 10856 70694
rect 1762 70632 1768 70644
rect 1596 70604 1768 70632
rect 1596 70573 1624 70604
rect 1762 70592 1768 70604
rect 1820 70592 1826 70644
rect 2406 70592 2412 70644
rect 2464 70632 2470 70644
rect 2501 70635 2559 70641
rect 2501 70632 2513 70635
rect 2464 70604 2513 70632
rect 2464 70592 2470 70604
rect 2501 70601 2513 70604
rect 2547 70601 2559 70635
rect 9953 70635 10011 70641
rect 9953 70632 9965 70635
rect 2501 70595 2559 70601
rect 6886 70604 9965 70632
rect 1581 70567 1639 70573
rect 1581 70533 1593 70567
rect 1627 70533 1639 70567
rect 1581 70527 1639 70533
rect 1673 70567 1731 70573
rect 1673 70533 1685 70567
rect 1719 70564 1731 70567
rect 6886 70564 6914 70604
rect 9953 70601 9965 70604
rect 9999 70601 10011 70635
rect 9953 70595 10011 70601
rect 1719 70536 6914 70564
rect 1719 70533 1731 70536
rect 1673 70527 1731 70533
rect 1302 70456 1308 70508
rect 1360 70496 1366 70508
rect 1397 70499 1455 70505
rect 1397 70496 1409 70499
rect 1360 70468 1409 70496
rect 1360 70456 1366 70468
rect 1397 70465 1409 70468
rect 1443 70465 1455 70499
rect 1397 70459 1455 70465
rect 1762 70456 1768 70508
rect 1820 70505 1826 70508
rect 1820 70496 1828 70505
rect 2590 70496 2596 70508
rect 1820 70468 2596 70496
rect 1820 70459 1828 70468
rect 1820 70456 1826 70459
rect 2590 70456 2596 70468
rect 2648 70456 2654 70508
rect 2685 70499 2743 70505
rect 2685 70465 2697 70499
rect 2731 70496 2743 70499
rect 2958 70496 2964 70508
rect 2731 70468 2964 70496
rect 2731 70465 2743 70468
rect 2685 70459 2743 70465
rect 2958 70456 2964 70468
rect 3016 70456 3022 70508
rect 10137 70499 10195 70505
rect 10137 70465 10149 70499
rect 10183 70465 10195 70499
rect 10137 70459 10195 70465
rect 5718 70428 5724 70440
rect 1964 70400 5724 70428
rect 1964 70369 1992 70400
rect 5718 70388 5724 70400
rect 5776 70388 5782 70440
rect 10152 70372 10180 70459
rect 1949 70363 2007 70369
rect 1949 70329 1961 70363
rect 1995 70360 2007 70363
rect 1995 70332 2029 70360
rect 1995 70329 2007 70332
rect 1949 70323 2007 70329
rect 10134 70320 10140 70372
rect 10192 70320 10198 70372
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5845 70202
rect 5897 70150 5909 70202
rect 5961 70150 5973 70202
rect 6025 70150 6037 70202
rect 6089 70150 6101 70202
rect 6153 70150 9109 70202
rect 9161 70150 9173 70202
rect 9225 70150 9237 70202
rect 9289 70150 9301 70202
rect 9353 70150 9365 70202
rect 9417 70150 10856 70202
rect 1104 70128 10856 70150
rect 1949 70023 2007 70029
rect 1949 69989 1961 70023
rect 1995 70020 2007 70023
rect 3602 70020 3608 70032
rect 1995 69992 3608 70020
rect 1995 69989 2007 69992
rect 1949 69983 2007 69989
rect 3602 69980 3608 69992
rect 3660 69980 3666 70032
rect 1394 69884 1400 69896
rect 1355 69856 1400 69884
rect 1394 69844 1400 69856
rect 1452 69844 1458 69896
rect 1578 69884 1584 69896
rect 1539 69856 1584 69884
rect 1578 69844 1584 69856
rect 1636 69844 1642 69896
rect 1762 69844 1768 69896
rect 1820 69893 1826 69896
rect 1820 69884 1828 69893
rect 2685 69887 2743 69893
rect 1820 69856 1865 69884
rect 1820 69847 1828 69856
rect 2685 69853 2697 69887
rect 2731 69884 2743 69887
rect 3050 69884 3056 69896
rect 2731 69856 3056 69884
rect 2731 69853 2743 69856
rect 2685 69847 2743 69853
rect 1820 69844 1826 69847
rect 3050 69844 3056 69856
rect 3108 69844 3114 69896
rect 10134 69884 10140 69896
rect 10095 69856 10140 69884
rect 10134 69844 10140 69856
rect 10192 69844 10198 69896
rect 1673 69819 1731 69825
rect 1673 69785 1685 69819
rect 1719 69816 1731 69819
rect 1719 69788 2774 69816
rect 1719 69785 1731 69788
rect 1673 69779 1731 69785
rect 1578 69708 1584 69760
rect 1636 69748 1642 69760
rect 2222 69748 2228 69760
rect 1636 69720 2228 69748
rect 1636 69708 1642 69720
rect 2222 69708 2228 69720
rect 2280 69708 2286 69760
rect 2501 69751 2559 69757
rect 2501 69717 2513 69751
rect 2547 69748 2559 69751
rect 2590 69748 2596 69760
rect 2547 69720 2596 69748
rect 2547 69717 2559 69720
rect 2501 69711 2559 69717
rect 2590 69708 2596 69720
rect 2648 69708 2654 69760
rect 2746 69748 2774 69788
rect 9953 69751 10011 69757
rect 9953 69748 9965 69751
rect 2746 69720 9965 69748
rect 9953 69717 9965 69720
rect 9999 69717 10011 69751
rect 9953 69711 10011 69717
rect 1104 69658 10856 69680
rect 1104 69606 4213 69658
rect 4265 69606 4277 69658
rect 4329 69606 4341 69658
rect 4393 69606 4405 69658
rect 4457 69606 4469 69658
rect 4521 69606 7477 69658
rect 7529 69606 7541 69658
rect 7593 69606 7605 69658
rect 7657 69606 7669 69658
rect 7721 69606 7733 69658
rect 7785 69606 10856 69658
rect 1104 69584 10856 69606
rect 1394 69504 1400 69556
rect 1452 69504 1458 69556
rect 1412 69417 1440 69504
rect 1581 69479 1639 69485
rect 1581 69445 1593 69479
rect 1627 69476 1639 69479
rect 1946 69476 1952 69488
rect 1627 69448 1952 69476
rect 1627 69445 1639 69448
rect 1581 69439 1639 69445
rect 1946 69436 1952 69448
rect 2004 69436 2010 69488
rect 1397 69411 1455 69417
rect 1397 69377 1409 69411
rect 1443 69377 1455 69411
rect 1397 69371 1455 69377
rect 1673 69411 1731 69417
rect 1673 69377 1685 69411
rect 1719 69377 1731 69411
rect 1673 69371 1731 69377
rect 1302 69300 1308 69352
rect 1360 69340 1366 69352
rect 1412 69340 1440 69371
rect 1360 69312 1440 69340
rect 1688 69340 1716 69371
rect 1762 69368 1768 69420
rect 1820 69417 1826 69420
rect 1820 69408 1828 69417
rect 2685 69411 2743 69417
rect 1820 69380 1865 69408
rect 1820 69371 1828 69380
rect 2685 69377 2697 69411
rect 2731 69408 2743 69411
rect 2958 69408 2964 69420
rect 2731 69380 2964 69408
rect 2731 69377 2743 69380
rect 2685 69371 2743 69377
rect 1820 69368 1826 69371
rect 2958 69368 2964 69380
rect 3016 69368 3022 69420
rect 3326 69408 3332 69420
rect 3287 69380 3332 69408
rect 3326 69368 3332 69380
rect 3384 69368 3390 69420
rect 9950 69340 9956 69352
rect 1688 69312 9956 69340
rect 1360 69300 1366 69312
rect 9950 69300 9956 69312
rect 10008 69300 10014 69352
rect 753 69275 811 69281
rect 753 69241 765 69275
rect 799 69272 811 69275
rect 2590 69272 2596 69284
rect 799 69244 2596 69272
rect 799 69241 811 69244
rect 753 69235 811 69241
rect 2590 69232 2596 69244
rect 2648 69232 2654 69284
rect 1210 69164 1216 69216
rect 1268 69204 1274 69216
rect 1949 69207 2007 69213
rect 1949 69204 1961 69207
rect 1268 69176 1961 69204
rect 1268 69164 1274 69176
rect 1949 69173 1961 69176
rect 1995 69173 2007 69207
rect 1949 69167 2007 69173
rect 2130 69164 2136 69216
rect 2188 69204 2194 69216
rect 2501 69207 2559 69213
rect 2501 69204 2513 69207
rect 2188 69176 2513 69204
rect 2188 69164 2194 69176
rect 2501 69173 2513 69176
rect 2547 69173 2559 69207
rect 2501 69167 2559 69173
rect 3145 69207 3203 69213
rect 3145 69173 3157 69207
rect 3191 69204 3203 69207
rect 3510 69204 3516 69216
rect 3191 69176 3516 69204
rect 3191 69173 3203 69176
rect 3145 69167 3203 69173
rect 3510 69164 3516 69176
rect 3568 69164 3574 69216
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5845 69114
rect 5897 69062 5909 69114
rect 5961 69062 5973 69114
rect 6025 69062 6037 69114
rect 6089 69062 6101 69114
rect 6153 69062 9109 69114
rect 9161 69062 9173 69114
rect 9225 69062 9237 69114
rect 9289 69062 9301 69114
rect 9353 69062 9365 69114
rect 9417 69062 10856 69114
rect 1104 69040 10856 69062
rect 1394 68960 1400 69012
rect 1452 69000 1458 69012
rect 1946 69000 1952 69012
rect 1452 68972 1952 69000
rect 1452 68960 1458 68972
rect 1946 68960 1952 68972
rect 2004 68960 2010 69012
rect 9950 69000 9956 69012
rect 9911 68972 9956 69000
rect 9950 68960 9956 68972
rect 10008 68960 10014 69012
rect 2590 68892 2596 68944
rect 2648 68892 2654 68944
rect 11057 68935 11115 68941
rect 11057 68932 11069 68935
rect 2700 68904 11069 68932
rect 1762 68824 1768 68876
rect 1820 68864 1826 68876
rect 2608 68864 2636 68892
rect 1820 68836 2636 68864
rect 1820 68824 1826 68836
rect 1394 68796 1400 68808
rect 1355 68768 1400 68796
rect 1394 68756 1400 68768
rect 1452 68756 1458 68808
rect 2511 68805 2539 68836
rect 2496 68799 2554 68805
rect 2496 68765 2508 68799
rect 2542 68765 2554 68799
rect 2496 68759 2554 68765
rect 2593 68799 2651 68805
rect 2593 68765 2605 68799
rect 2639 68796 2651 68799
rect 2700 68796 2728 68904
rect 11057 68901 11069 68904
rect 11103 68901 11115 68935
rect 11057 68895 11115 68901
rect 2866 68796 2872 68808
rect 2639 68768 2728 68796
rect 2827 68768 2872 68796
rect 2639 68765 2651 68768
rect 2593 68759 2651 68765
rect 2866 68756 2872 68768
rect 2924 68756 2930 68808
rect 10134 68796 10140 68808
rect 10095 68768 10140 68796
rect 10134 68756 10140 68768
rect 10192 68756 10198 68808
rect 2685 68731 2743 68737
rect 2685 68697 2697 68731
rect 2731 68728 2743 68731
rect 3418 68728 3424 68740
rect 2731 68700 3424 68728
rect 2731 68697 2743 68700
rect 2685 68691 2743 68697
rect 3418 68688 3424 68700
rect 3476 68688 3482 68740
rect 1581 68663 1639 68669
rect 1581 68629 1593 68663
rect 1627 68660 1639 68663
rect 1762 68660 1768 68672
rect 1627 68632 1768 68660
rect 1627 68629 1639 68632
rect 1581 68623 1639 68629
rect 1762 68620 1768 68632
rect 1820 68620 1826 68672
rect 2309 68663 2367 68669
rect 2309 68629 2321 68663
rect 2355 68660 2367 68663
rect 7006 68660 7012 68672
rect 2355 68632 7012 68660
rect 2355 68629 2367 68632
rect 2309 68623 2367 68629
rect 7006 68620 7012 68632
rect 7064 68620 7070 68672
rect 1104 68570 10856 68592
rect 1104 68518 4213 68570
rect 4265 68518 4277 68570
rect 4329 68518 4341 68570
rect 4393 68518 4405 68570
rect 4457 68518 4469 68570
rect 4521 68518 7477 68570
rect 7529 68518 7541 68570
rect 7593 68518 7605 68570
rect 7657 68518 7669 68570
rect 7721 68518 7733 68570
rect 7785 68518 10856 68570
rect 1104 68496 10856 68518
rect 1578 68416 1584 68468
rect 1636 68416 1642 68468
rect 9953 68459 10011 68465
rect 9953 68456 9965 68459
rect 2976 68428 9965 68456
rect 1596 68388 1624 68416
rect 1596 68360 1808 68388
rect 1026 68280 1032 68332
rect 1084 68320 1090 68332
rect 1673 68323 1731 68329
rect 1673 68320 1685 68323
rect 1084 68292 1685 68320
rect 1084 68280 1090 68292
rect 1673 68289 1685 68292
rect 1719 68289 1731 68323
rect 1673 68283 1731 68289
rect 1302 68212 1308 68264
rect 1360 68252 1366 68264
rect 1397 68255 1455 68261
rect 1397 68252 1409 68255
rect 1360 68224 1409 68252
rect 1360 68212 1366 68224
rect 1397 68221 1409 68224
rect 1443 68221 1455 68255
rect 1397 68215 1455 68221
rect 1670 68144 1676 68196
rect 1728 68184 1734 68196
rect 1780 68184 1808 68360
rect 1946 68348 1952 68400
rect 2004 68388 2010 68400
rect 2976 68397 3004 68428
rect 9953 68425 9965 68428
rect 9999 68425 10011 68459
rect 9953 68419 10011 68425
rect 2869 68391 2927 68397
rect 2869 68388 2881 68391
rect 2004 68360 2881 68388
rect 2004 68348 2010 68360
rect 2869 68357 2881 68360
rect 2915 68357 2927 68391
rect 2869 68351 2927 68357
rect 2961 68391 3019 68397
rect 2961 68357 2973 68391
rect 3007 68357 3019 68391
rect 2961 68351 3019 68357
rect 2685 68323 2743 68329
rect 2685 68289 2697 68323
rect 2731 68320 2743 68323
rect 2774 68320 2780 68332
rect 2731 68292 2780 68320
rect 2731 68289 2743 68292
rect 2685 68283 2743 68289
rect 2774 68280 2780 68292
rect 2832 68280 2838 68332
rect 3050 68280 3056 68332
rect 3108 68329 3114 68332
rect 3108 68320 3116 68329
rect 10134 68320 10140 68332
rect 3108 68292 3153 68320
rect 10095 68292 10140 68320
rect 3108 68283 3116 68292
rect 3108 68280 3114 68283
rect 10134 68280 10140 68292
rect 10192 68280 10198 68332
rect 2590 68212 2596 68264
rect 2648 68252 2654 68264
rect 3068 68252 3096 68280
rect 2648 68224 3096 68252
rect 2648 68212 2654 68224
rect 1728 68156 1808 68184
rect 1728 68144 1734 68156
rect 3237 68119 3295 68125
rect 3237 68085 3249 68119
rect 3283 68116 3295 68119
rect 5166 68116 5172 68128
rect 3283 68088 5172 68116
rect 3283 68085 3295 68088
rect 3237 68079 3295 68085
rect 5166 68076 5172 68088
rect 5224 68076 5230 68128
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5845 68026
rect 5897 67974 5909 68026
rect 5961 67974 5973 68026
rect 6025 67974 6037 68026
rect 6089 67974 6101 68026
rect 6153 67974 9109 68026
rect 9161 67974 9173 68026
rect 9225 67974 9237 68026
rect 9289 67974 9301 68026
rect 9353 67974 9365 68026
rect 9417 67974 10856 68026
rect 1104 67952 10856 67974
rect 1118 67736 1124 67788
rect 1176 67776 1182 67788
rect 1673 67779 1731 67785
rect 1673 67776 1685 67779
rect 1176 67748 1685 67776
rect 1176 67736 1182 67748
rect 1673 67745 1685 67748
rect 1719 67745 1731 67779
rect 1673 67739 1731 67745
rect 1394 67708 1400 67720
rect 1355 67680 1400 67708
rect 1394 67668 1400 67680
rect 1452 67668 1458 67720
rect 1104 67482 10856 67504
rect 1104 67430 4213 67482
rect 4265 67430 4277 67482
rect 4329 67430 4341 67482
rect 4393 67430 4405 67482
rect 4457 67430 4469 67482
rect 4521 67430 7477 67482
rect 7529 67430 7541 67482
rect 7593 67430 7605 67482
rect 7657 67430 7669 67482
rect 7721 67430 7733 67482
rect 7785 67430 10856 67482
rect 1104 67408 10856 67430
rect 382 67192 388 67244
rect 440 67232 446 67244
rect 1673 67235 1731 67241
rect 1673 67232 1685 67235
rect 440 67204 1685 67232
rect 440 67192 446 67204
rect 1673 67201 1685 67204
rect 1719 67201 1731 67235
rect 10134 67232 10140 67244
rect 10095 67204 10140 67232
rect 1673 67195 1731 67201
rect 10134 67192 10140 67204
rect 10192 67192 10198 67244
rect 1394 67164 1400 67176
rect 1355 67136 1400 67164
rect 1394 67124 1400 67136
rect 1452 67124 1458 67176
rect 9950 67028 9956 67040
rect 9911 67000 9956 67028
rect 9950 66988 9956 67000
rect 10008 66988 10014 67040
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5845 66938
rect 5897 66886 5909 66938
rect 5961 66886 5973 66938
rect 6025 66886 6037 66938
rect 6089 66886 6101 66938
rect 6153 66886 9109 66938
rect 9161 66886 9173 66938
rect 9225 66886 9237 66938
rect 9289 66886 9301 66938
rect 9353 66886 9365 66938
rect 9417 66886 10856 66938
rect 1104 66864 10856 66886
rect 3234 66716 3240 66768
rect 3292 66756 3298 66768
rect 3786 66756 3792 66768
rect 3292 66728 3792 66756
rect 3292 66716 3298 66728
rect 3786 66716 3792 66728
rect 3844 66716 3850 66768
rect 1394 66620 1400 66632
rect 1355 66592 1400 66620
rect 1394 66580 1400 66592
rect 1452 66580 1458 66632
rect 1673 66623 1731 66629
rect 1673 66589 1685 66623
rect 1719 66620 1731 66623
rect 1854 66620 1860 66632
rect 1719 66592 1860 66620
rect 1719 66589 1731 66592
rect 1673 66583 1731 66589
rect 1854 66580 1860 66592
rect 1912 66580 1918 66632
rect 2961 66623 3019 66629
rect 2961 66589 2973 66623
rect 3007 66620 3019 66623
rect 3234 66620 3240 66632
rect 3007 66592 3240 66620
rect 3007 66589 3019 66592
rect 2961 66583 3019 66589
rect 3234 66580 3240 66592
rect 3292 66580 3298 66632
rect 10134 66620 10140 66632
rect 10095 66592 10140 66620
rect 10134 66580 10140 66592
rect 10192 66580 10198 66632
rect 2314 66512 2320 66564
rect 2372 66552 2378 66564
rect 3142 66552 3148 66564
rect 2372 66524 3148 66552
rect 2372 66512 2378 66524
rect 3142 66512 3148 66524
rect 3200 66512 3206 66564
rect 845 66487 903 66493
rect 845 66453 857 66487
rect 891 66484 903 66487
rect 2222 66484 2228 66496
rect 891 66456 2228 66484
rect 891 66453 903 66456
rect 845 66447 903 66453
rect 2222 66444 2228 66456
rect 2280 66444 2286 66496
rect 2777 66487 2835 66493
rect 2777 66453 2789 66487
rect 2823 66484 2835 66487
rect 2958 66484 2964 66496
rect 2823 66456 2964 66484
rect 2823 66453 2835 66456
rect 2777 66447 2835 66453
rect 2958 66444 2964 66456
rect 3016 66444 3022 66496
rect 9858 66444 9864 66496
rect 9916 66484 9922 66496
rect 9953 66487 10011 66493
rect 9953 66484 9965 66487
rect 9916 66456 9965 66484
rect 9916 66444 9922 66456
rect 9953 66453 9965 66456
rect 9999 66453 10011 66487
rect 9953 66447 10011 66453
rect 1104 66394 10856 66416
rect 1104 66342 4213 66394
rect 4265 66342 4277 66394
rect 4329 66342 4341 66394
rect 4393 66342 4405 66394
rect 4457 66342 4469 66394
rect 4521 66342 7477 66394
rect 7529 66342 7541 66394
rect 7593 66342 7605 66394
rect 7657 66342 7669 66394
rect 7721 66342 7733 66394
rect 7785 66342 10856 66394
rect 1104 66320 10856 66342
rect 1302 66240 1308 66292
rect 1360 66280 1366 66292
rect 1670 66280 1676 66292
rect 1360 66252 1676 66280
rect 1360 66240 1366 66252
rect 1670 66240 1676 66252
rect 1728 66240 1734 66292
rect 2866 66280 2872 66292
rect 1872 66252 2355 66280
rect 1578 66212 1584 66224
rect 1539 66184 1584 66212
rect 1578 66172 1584 66184
rect 1636 66172 1642 66224
rect 1872 66212 1900 66252
rect 1832 66184 1900 66212
rect 937 66147 995 66153
rect 937 66113 949 66147
rect 983 66144 995 66147
rect 1397 66147 1455 66153
rect 1397 66144 1409 66147
rect 983 66116 1409 66144
rect 983 66113 995 66116
rect 937 66107 995 66113
rect 1397 66113 1409 66116
rect 1443 66113 1455 66147
rect 1670 66144 1676 66156
rect 1631 66116 1676 66144
rect 1397 66107 1455 66113
rect 1670 66104 1676 66116
rect 1728 66104 1734 66156
rect 1832 66153 1860 66184
rect 1817 66147 1875 66153
rect 1817 66113 1829 66147
rect 1863 66113 1875 66147
rect 1817 66107 1875 66113
rect 2222 66036 2228 66088
rect 2280 66076 2286 66088
rect 2327 66076 2355 66252
rect 2516 66252 2872 66280
rect 2516 66156 2544 66252
rect 2866 66240 2872 66252
rect 2924 66240 2930 66292
rect 2590 66172 2596 66224
rect 2648 66212 2654 66224
rect 2685 66215 2743 66221
rect 2685 66212 2697 66215
rect 2648 66184 2697 66212
rect 2648 66172 2654 66184
rect 2685 66181 2697 66184
rect 2731 66181 2743 66215
rect 2685 66175 2743 66181
rect 2777 66215 2835 66221
rect 2777 66181 2789 66215
rect 2823 66212 2835 66215
rect 9950 66212 9956 66224
rect 2823 66184 9956 66212
rect 2823 66181 2835 66184
rect 2777 66175 2835 66181
rect 9950 66172 9956 66184
rect 10008 66172 10014 66224
rect 2498 66144 2504 66156
rect 2459 66116 2504 66144
rect 2498 66104 2504 66116
rect 2556 66104 2562 66156
rect 2921 66147 2979 66153
rect 2921 66113 2933 66147
rect 2967 66144 2979 66147
rect 3050 66144 3056 66156
rect 2967 66116 3056 66144
rect 2967 66113 2979 66116
rect 2921 66107 2979 66113
rect 3050 66104 3056 66116
rect 3108 66104 3114 66156
rect 10134 66144 10140 66156
rect 10095 66116 10140 66144
rect 10134 66104 10140 66116
rect 10192 66104 10198 66156
rect 2280 66048 2355 66076
rect 2280 66036 2286 66048
rect 1949 66011 2007 66017
rect 1949 65977 1961 66011
rect 1995 66008 2007 66011
rect 7098 66008 7104 66020
rect 1995 65980 7104 66008
rect 1995 65977 2007 65980
rect 1949 65971 2007 65977
rect 7098 65968 7104 65980
rect 7156 65968 7162 66020
rect 7190 65968 7196 66020
rect 7248 66008 7254 66020
rect 9953 66011 10011 66017
rect 9953 66008 9965 66011
rect 7248 65980 9965 66008
rect 7248 65968 7254 65980
rect 9953 65977 9965 65980
rect 9999 65977 10011 66011
rect 9953 65971 10011 65977
rect 3053 65943 3111 65949
rect 3053 65909 3065 65943
rect 3099 65940 3111 65943
rect 11425 65943 11483 65949
rect 11425 65940 11437 65943
rect 3099 65912 11437 65940
rect 3099 65909 3111 65912
rect 3053 65903 3111 65909
rect 11425 65909 11437 65912
rect 11471 65909 11483 65943
rect 11425 65903 11483 65909
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5845 65850
rect 5897 65798 5909 65850
rect 5961 65798 5973 65850
rect 6025 65798 6037 65850
rect 6089 65798 6101 65850
rect 6153 65798 9109 65850
rect 9161 65798 9173 65850
rect 9225 65798 9237 65850
rect 9289 65798 9301 65850
rect 9353 65798 9365 65850
rect 9417 65798 10856 65850
rect 1104 65776 10856 65798
rect 11241 65807 11299 65813
rect 11241 65773 11253 65807
rect 11287 65804 11299 65807
rect 11609 65807 11667 65813
rect 11609 65804 11621 65807
rect 11287 65776 11621 65804
rect 11287 65773 11299 65776
rect 11241 65767 11299 65773
rect 11609 65773 11621 65776
rect 11655 65773 11667 65807
rect 11609 65767 11667 65773
rect 2424 65708 5396 65736
rect 1762 65628 1768 65680
rect 1820 65668 1826 65680
rect 2133 65671 2191 65677
rect 2133 65668 2145 65671
rect 1820 65640 2145 65668
rect 1820 65628 1826 65640
rect 2133 65637 2145 65640
rect 2179 65637 2191 65671
rect 2133 65631 2191 65637
rect 1670 65560 1676 65612
rect 1728 65600 1734 65612
rect 1946 65600 1952 65612
rect 1728 65572 1952 65600
rect 1728 65560 1734 65572
rect 1946 65560 1952 65572
rect 2004 65560 2010 65612
rect 1394 65532 1400 65544
rect 1355 65504 1400 65532
rect 1394 65492 1400 65504
rect 1452 65492 1458 65544
rect 2424 65541 2452 65708
rect 3142 65668 3148 65680
rect 2521 65640 3148 65668
rect 2521 65541 2549 65640
rect 3142 65628 3148 65640
rect 3200 65628 3206 65680
rect 5368 65600 5396 65708
rect 7098 65696 7104 65748
rect 7156 65736 7162 65748
rect 11333 65739 11391 65745
rect 11333 65736 11345 65739
rect 7156 65708 11345 65736
rect 7156 65696 7162 65708
rect 11333 65705 11345 65708
rect 11379 65705 11391 65739
rect 11333 65699 11391 65705
rect 5902 65628 5908 65680
rect 5960 65668 5966 65680
rect 11241 65671 11299 65677
rect 11241 65668 11253 65671
rect 5960 65640 11253 65668
rect 5960 65628 5966 65640
rect 11241 65637 11253 65640
rect 11287 65637 11299 65671
rect 11241 65631 11299 65637
rect 9858 65600 9864 65612
rect 5368 65572 9864 65600
rect 9858 65560 9864 65572
rect 9916 65560 9922 65612
rect 2265 65535 2323 65541
rect 2265 65532 2277 65535
rect 2240 65501 2277 65532
rect 2311 65501 2323 65535
rect 2240 65495 2323 65501
rect 2409 65535 2467 65541
rect 2409 65501 2421 65535
rect 2455 65501 2467 65535
rect 2521 65535 2605 65541
rect 2521 65504 2559 65535
rect 2409 65495 2467 65501
rect 2547 65501 2559 65504
rect 2593 65501 2605 65535
rect 2547 65495 2605 65501
rect 2240 65464 2268 65495
rect 2682 65492 2688 65544
rect 2740 65532 2746 65544
rect 3789 65535 3847 65541
rect 2740 65504 2785 65532
rect 2740 65492 2746 65504
rect 3789 65501 3801 65535
rect 3835 65501 3847 65535
rect 3789 65495 3847 65501
rect 3050 65464 3056 65476
rect 2240 65436 3056 65464
rect 3050 65424 3056 65436
rect 3108 65424 3114 65476
rect 3142 65424 3148 65476
rect 3200 65464 3206 65476
rect 3804 65464 3832 65495
rect 3200 65436 3832 65464
rect 3200 65424 3206 65436
rect 1581 65399 1639 65405
rect 1581 65365 1593 65399
rect 1627 65396 1639 65399
rect 1762 65396 1768 65408
rect 1627 65368 1768 65396
rect 1627 65365 1639 65368
rect 1581 65359 1639 65365
rect 1762 65356 1768 65368
rect 1820 65356 1826 65408
rect 3326 65356 3332 65408
rect 3384 65396 3390 65408
rect 3973 65399 4031 65405
rect 3973 65396 3985 65399
rect 3384 65368 3985 65396
rect 3384 65356 3390 65368
rect 3973 65365 3985 65368
rect 4019 65365 4031 65399
rect 3973 65359 4031 65365
rect 1104 65306 10856 65328
rect 1104 65254 4213 65306
rect 4265 65254 4277 65306
rect 4329 65254 4341 65306
rect 4393 65254 4405 65306
rect 4457 65254 4469 65306
rect 4521 65254 7477 65306
rect 7529 65254 7541 65306
rect 7593 65254 7605 65306
rect 7657 65254 7669 65306
rect 7721 65254 7733 65306
rect 7785 65254 10856 65306
rect 1104 65232 10856 65254
rect 1949 65195 2007 65201
rect 1949 65161 1961 65195
rect 1995 65192 2007 65195
rect 6822 65192 6828 65204
rect 1995 65164 6828 65192
rect 1995 65161 2007 65164
rect 1949 65155 2007 65161
rect 6822 65152 6828 65164
rect 6880 65152 6886 65204
rect 845 65127 903 65133
rect 845 65093 857 65127
rect 891 65124 903 65127
rect 1581 65127 1639 65133
rect 1581 65124 1593 65127
rect 891 65096 1593 65124
rect 891 65093 903 65096
rect 845 65087 903 65093
rect 1581 65093 1593 65096
rect 1627 65093 1639 65127
rect 1581 65087 1639 65093
rect 1673 65127 1731 65133
rect 1673 65093 1685 65127
rect 1719 65124 1731 65127
rect 11517 65127 11575 65133
rect 11517 65124 11529 65127
rect 1719 65096 11529 65124
rect 1719 65093 1731 65096
rect 1673 65087 1731 65093
rect 11517 65093 11529 65096
rect 11563 65093 11575 65127
rect 11517 65087 11575 65093
rect 937 65059 995 65065
rect 937 65025 949 65059
rect 983 65056 995 65059
rect 1397 65059 1455 65065
rect 1397 65056 1409 65059
rect 983 65028 1409 65056
rect 983 65025 995 65028
rect 937 65019 995 65025
rect 1397 65025 1409 65028
rect 1443 65025 1455 65059
rect 1397 65019 1455 65025
rect 1765 65059 1823 65065
rect 1765 65025 1777 65059
rect 1811 65056 1823 65059
rect 2038 65056 2044 65068
rect 1811 65028 2044 65056
rect 1811 65025 1823 65028
rect 1765 65019 1823 65025
rect 2038 65016 2044 65028
rect 2096 65056 2102 65068
rect 2222 65056 2228 65068
rect 2096 65028 2228 65056
rect 2096 65016 2102 65028
rect 2222 65016 2228 65028
rect 2280 65016 2286 65068
rect 2961 65059 3019 65065
rect 2961 65025 2973 65059
rect 3007 65056 3019 65059
rect 3050 65056 3056 65068
rect 3007 65028 3056 65056
rect 3007 65025 3019 65028
rect 2961 65019 3019 65025
rect 3050 65016 3056 65028
rect 3108 65016 3114 65068
rect 3237 65059 3295 65065
rect 3237 65025 3249 65059
rect 3283 65056 3295 65059
rect 3418 65056 3424 65068
rect 3283 65028 3424 65056
rect 3283 65025 3295 65028
rect 3237 65019 3295 65025
rect 3418 65016 3424 65028
rect 3476 65016 3482 65068
rect 3697 65059 3755 65065
rect 3697 65025 3709 65059
rect 3743 65025 3755 65059
rect 10134 65056 10140 65068
rect 10095 65028 10140 65056
rect 3697 65019 3755 65025
rect 3712 64988 3740 65019
rect 10134 65016 10140 65028
rect 10192 65016 10198 65068
rect 2148 64960 3740 64988
rect 2148 64864 2176 64960
rect 3878 64920 3884 64932
rect 3839 64892 3884 64920
rect 3878 64880 3884 64892
rect 3936 64880 3942 64932
rect 2130 64812 2136 64864
rect 2188 64812 2194 64864
rect 3418 64812 3424 64864
rect 3476 64852 3482 64864
rect 3602 64852 3608 64864
rect 3476 64824 3608 64852
rect 3476 64812 3482 64824
rect 3602 64812 3608 64824
rect 3660 64812 3666 64864
rect 6362 64812 6368 64864
rect 6420 64852 6426 64864
rect 9953 64855 10011 64861
rect 9953 64852 9965 64855
rect 6420 64824 9965 64852
rect 6420 64812 6426 64824
rect 9953 64821 9965 64824
rect 9999 64821 10011 64855
rect 9953 64815 10011 64821
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5845 64762
rect 5897 64710 5909 64762
rect 5961 64710 5973 64762
rect 6025 64710 6037 64762
rect 6089 64710 6101 64762
rect 6153 64710 9109 64762
rect 9161 64710 9173 64762
rect 9225 64710 9237 64762
rect 9289 64710 9301 64762
rect 9353 64710 9365 64762
rect 9417 64710 10856 64762
rect 1104 64688 10856 64710
rect 1949 64583 2007 64589
rect 1949 64549 1961 64583
rect 1995 64580 2007 64583
rect 6914 64580 6920 64592
rect 1995 64552 6920 64580
rect 1995 64549 2007 64552
rect 1949 64543 2007 64549
rect 6914 64540 6920 64552
rect 6972 64540 6978 64592
rect 937 64447 995 64453
rect 937 64413 949 64447
rect 983 64444 995 64447
rect 1397 64447 1455 64453
rect 1397 64444 1409 64447
rect 983 64416 1409 64444
rect 983 64413 995 64416
rect 937 64407 995 64413
rect 1397 64413 1409 64416
rect 1443 64413 1455 64447
rect 1397 64407 1455 64413
rect 1486 64404 1492 64456
rect 1544 64444 1550 64456
rect 1581 64447 1639 64453
rect 1581 64444 1593 64447
rect 1544 64416 1593 64444
rect 1544 64404 1550 64416
rect 1581 64413 1593 64416
rect 1627 64413 1639 64447
rect 1581 64407 1639 64413
rect 1817 64447 1875 64453
rect 1817 64413 1829 64447
rect 1863 64444 1875 64447
rect 2038 64444 2044 64456
rect 1863 64416 2044 64444
rect 1863 64413 1875 64416
rect 1817 64407 1875 64413
rect 2038 64404 2044 64416
rect 2096 64404 2102 64456
rect 2222 64404 2228 64456
rect 2280 64444 2286 64456
rect 2501 64447 2559 64453
rect 2501 64444 2513 64447
rect 2280 64416 2513 64444
rect 2280 64404 2286 64416
rect 2501 64413 2513 64416
rect 2547 64413 2559 64447
rect 10134 64444 10140 64456
rect 10095 64416 10140 64444
rect 2501 64407 2559 64413
rect 10134 64404 10140 64416
rect 10192 64404 10198 64456
rect 1673 64379 1731 64385
rect 1673 64345 1685 64379
rect 1719 64376 1731 64379
rect 6362 64376 6368 64388
rect 1719 64348 6368 64376
rect 1719 64345 1731 64348
rect 1673 64339 1731 64345
rect 6362 64336 6368 64348
rect 6420 64336 6426 64388
rect 2685 64311 2743 64317
rect 2685 64277 2697 64311
rect 2731 64308 2743 64311
rect 2774 64308 2780 64320
rect 2731 64280 2780 64308
rect 2731 64277 2743 64280
rect 2685 64271 2743 64277
rect 2774 64268 2780 64280
rect 2832 64268 2838 64320
rect 9950 64308 9956 64320
rect 9911 64280 9956 64308
rect 9950 64268 9956 64280
rect 10008 64268 10014 64320
rect 1104 64218 10856 64240
rect 1104 64166 4213 64218
rect 4265 64166 4277 64218
rect 4329 64166 4341 64218
rect 4393 64166 4405 64218
rect 4457 64166 4469 64218
rect 4521 64166 7477 64218
rect 7529 64166 7541 64218
rect 7593 64166 7605 64218
rect 7657 64166 7669 64218
rect 7721 64166 7733 64218
rect 7785 64166 10856 64218
rect 1104 64144 10856 64166
rect 937 64039 995 64045
rect 937 64005 949 64039
rect 983 64036 995 64039
rect 2222 64036 2228 64048
rect 983 64008 2228 64036
rect 983 64005 995 64008
rect 937 63999 995 64005
rect 2222 63996 2228 64008
rect 2280 63996 2286 64048
rect 1673 63971 1731 63977
rect 1673 63937 1685 63971
rect 1719 63937 1731 63971
rect 1673 63931 1731 63937
rect 2409 63971 2467 63977
rect 2409 63937 2421 63971
rect 2455 63968 2467 63971
rect 3694 63968 3700 63980
rect 2455 63940 3700 63968
rect 2455 63937 2467 63940
rect 2409 63931 2467 63937
rect 1688 63900 1716 63931
rect 3694 63928 3700 63940
rect 3752 63928 3758 63980
rect 4614 63900 4620 63912
rect 1688 63872 4620 63900
rect 4614 63860 4620 63872
rect 4672 63860 4678 63912
rect 1394 63724 1400 63776
rect 1452 63764 1458 63776
rect 1489 63767 1547 63773
rect 1489 63764 1501 63767
rect 1452 63736 1501 63764
rect 1452 63724 1458 63736
rect 1489 63733 1501 63736
rect 1535 63733 1547 63767
rect 2222 63764 2228 63776
rect 2183 63736 2228 63764
rect 1489 63727 1547 63733
rect 2222 63724 2228 63736
rect 2280 63724 2286 63776
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5845 63674
rect 5897 63622 5909 63674
rect 5961 63622 5973 63674
rect 6025 63622 6037 63674
rect 6089 63622 6101 63674
rect 6153 63622 9109 63674
rect 9161 63622 9173 63674
rect 9225 63622 9237 63674
rect 9289 63622 9301 63674
rect 9353 63622 9365 63674
rect 9417 63622 10856 63674
rect 1104 63600 10856 63622
rect 2317 63495 2375 63501
rect 2317 63461 2329 63495
rect 2363 63492 2375 63495
rect 2866 63492 2872 63504
rect 2363 63464 2872 63492
rect 2363 63461 2375 63464
rect 2317 63455 2375 63461
rect 2866 63452 2872 63464
rect 2924 63452 2930 63504
rect 934 63316 940 63368
rect 992 63356 998 63368
rect 1673 63359 1731 63365
rect 1673 63356 1685 63359
rect 992 63328 1685 63356
rect 992 63316 998 63328
rect 1673 63325 1685 63328
rect 1719 63325 1731 63359
rect 1673 63319 1731 63325
rect 2038 63316 2044 63368
rect 2096 63356 2102 63368
rect 2133 63359 2191 63365
rect 2133 63356 2145 63359
rect 2096 63328 2145 63356
rect 2096 63316 2102 63328
rect 2133 63325 2145 63328
rect 2179 63325 2191 63359
rect 2133 63319 2191 63325
rect 2498 63316 2504 63368
rect 2556 63356 2562 63368
rect 2869 63359 2927 63365
rect 2869 63356 2881 63359
rect 2556 63328 2881 63356
rect 2556 63316 2562 63328
rect 2869 63325 2881 63328
rect 2915 63325 2927 63359
rect 10134 63356 10140 63368
rect 10095 63328 10140 63356
rect 2869 63319 2927 63325
rect 10134 63316 10140 63328
rect 10192 63316 10198 63368
rect 1486 63220 1492 63232
rect 1447 63192 1492 63220
rect 1486 63180 1492 63192
rect 1544 63180 1550 63232
rect 3050 63220 3056 63232
rect 3011 63192 3056 63220
rect 3050 63180 3056 63192
rect 3108 63180 3114 63232
rect 9858 63180 9864 63232
rect 9916 63220 9922 63232
rect 9953 63223 10011 63229
rect 9953 63220 9965 63223
rect 9916 63192 9965 63220
rect 9916 63180 9922 63192
rect 9953 63189 9965 63192
rect 9999 63189 10011 63223
rect 9953 63183 10011 63189
rect 1104 63130 10856 63152
rect 1104 63078 4213 63130
rect 4265 63078 4277 63130
rect 4329 63078 4341 63130
rect 4393 63078 4405 63130
rect 4457 63078 4469 63130
rect 4521 63078 7477 63130
rect 7529 63078 7541 63130
rect 7593 63078 7605 63130
rect 7657 63078 7669 63130
rect 7721 63078 7733 63130
rect 7785 63078 10856 63130
rect 1104 63056 10856 63078
rect 1578 62948 1584 62960
rect 1539 62920 1584 62948
rect 1578 62908 1584 62920
rect 1636 62908 1642 62960
rect 1673 62951 1731 62957
rect 1673 62917 1685 62951
rect 1719 62948 1731 62951
rect 9950 62948 9956 62960
rect 1719 62920 9956 62948
rect 1719 62917 1731 62920
rect 1673 62911 1731 62917
rect 9950 62908 9956 62920
rect 10008 62908 10014 62960
rect 845 62883 903 62889
rect 845 62849 857 62883
rect 891 62880 903 62883
rect 1397 62883 1455 62889
rect 1397 62880 1409 62883
rect 891 62852 1409 62880
rect 891 62849 903 62852
rect 845 62843 903 62849
rect 1397 62849 1409 62852
rect 1443 62849 1455 62883
rect 1397 62843 1455 62849
rect 1817 62883 1875 62889
rect 1817 62849 1829 62883
rect 1863 62880 1875 62883
rect 2130 62880 2136 62892
rect 1863 62852 2136 62880
rect 1863 62849 1875 62852
rect 1817 62843 1875 62849
rect 2130 62840 2136 62852
rect 2188 62880 2194 62892
rect 2869 62883 2927 62889
rect 2869 62880 2881 62883
rect 2188 62852 2881 62880
rect 2188 62840 2194 62852
rect 2869 62849 2881 62852
rect 2915 62849 2927 62883
rect 2869 62843 2927 62849
rect 3145 62883 3203 62889
rect 3145 62849 3157 62883
rect 3191 62880 3203 62883
rect 3326 62880 3332 62892
rect 3191 62852 3332 62880
rect 3191 62849 3203 62852
rect 3145 62843 3203 62849
rect 3326 62840 3332 62852
rect 3384 62840 3390 62892
rect 10134 62880 10140 62892
rect 10095 62852 10140 62880
rect 10134 62840 10140 62852
rect 10192 62840 10198 62892
rect 1949 62747 2007 62753
rect 1949 62713 1961 62747
rect 1995 62744 2007 62747
rect 8478 62744 8484 62756
rect 1995 62716 8484 62744
rect 1995 62713 2007 62716
rect 1949 62707 2007 62713
rect 8478 62704 8484 62716
rect 8536 62704 8542 62756
rect 9953 62679 10011 62685
rect 9953 62645 9965 62679
rect 9999 62676 10011 62679
rect 11057 62679 11115 62685
rect 11057 62676 11069 62679
rect 9999 62648 11069 62676
rect 9999 62645 10011 62648
rect 9953 62639 10011 62645
rect 11057 62645 11069 62648
rect 11103 62645 11115 62679
rect 11057 62639 11115 62645
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5845 62586
rect 5897 62534 5909 62586
rect 5961 62534 5973 62586
rect 6025 62534 6037 62586
rect 6089 62534 6101 62586
rect 6153 62534 9109 62586
rect 9161 62534 9173 62586
rect 9225 62534 9237 62586
rect 9289 62534 9301 62586
rect 9353 62534 9365 62586
rect 9417 62534 10856 62586
rect 1104 62512 10856 62534
rect 1394 62296 1400 62348
rect 1452 62336 1458 62348
rect 2038 62336 2044 62348
rect 1452 62308 2044 62336
rect 1452 62296 1458 62308
rect 2038 62296 2044 62308
rect 2096 62296 2102 62348
rect 2406 62296 2412 62348
rect 2464 62336 2470 62348
rect 2685 62339 2743 62345
rect 2685 62336 2697 62339
rect 2464 62308 2697 62336
rect 2464 62296 2470 62308
rect 2685 62305 2697 62308
rect 2731 62305 2743 62339
rect 2685 62299 2743 62305
rect 842 62228 848 62280
rect 900 62268 906 62280
rect 1673 62271 1731 62277
rect 1673 62268 1685 62271
rect 900 62240 1685 62268
rect 900 62228 906 62240
rect 1673 62237 1685 62240
rect 1719 62237 1731 62271
rect 2958 62268 2964 62280
rect 2919 62240 2964 62268
rect 1673 62231 1731 62237
rect 2958 62228 2964 62240
rect 3016 62228 3022 62280
rect 10134 62268 10140 62280
rect 10095 62240 10140 62268
rect 10134 62228 10140 62240
rect 10192 62228 10198 62280
rect 1394 62092 1400 62144
rect 1452 62132 1458 62144
rect 1489 62135 1547 62141
rect 1489 62132 1501 62135
rect 1452 62104 1501 62132
rect 1452 62092 1458 62104
rect 1489 62101 1501 62104
rect 1535 62101 1547 62135
rect 1489 62095 1547 62101
rect 9766 62092 9772 62144
rect 9824 62132 9830 62144
rect 9953 62135 10011 62141
rect 9953 62132 9965 62135
rect 9824 62104 9965 62132
rect 9824 62092 9830 62104
rect 9953 62101 9965 62104
rect 9999 62101 10011 62135
rect 9953 62095 10011 62101
rect 1104 62042 10856 62064
rect 1104 61990 4213 62042
rect 4265 61990 4277 62042
rect 4329 61990 4341 62042
rect 4393 61990 4405 62042
rect 4457 61990 4469 62042
rect 4521 61990 7477 62042
rect 7529 61990 7541 62042
rect 7593 61990 7605 62042
rect 7657 61990 7669 62042
rect 7721 61990 7733 62042
rect 7785 61990 10856 62042
rect 1104 61968 10856 61990
rect 198 61752 204 61804
rect 256 61792 262 61804
rect 1673 61795 1731 61801
rect 1673 61792 1685 61795
rect 256 61764 1685 61792
rect 256 61752 262 61764
rect 1673 61761 1685 61764
rect 1719 61761 1731 61795
rect 1673 61755 1731 61761
rect 2038 61752 2044 61804
rect 2096 61792 2102 61804
rect 2409 61795 2467 61801
rect 2409 61792 2421 61795
rect 2096 61764 2421 61792
rect 2096 61752 2102 61764
rect 2409 61761 2421 61764
rect 2455 61761 2467 61795
rect 2409 61755 2467 61761
rect 1486 61684 1492 61736
rect 1544 61724 1550 61736
rect 1544 61696 2268 61724
rect 1544 61684 1550 61696
rect 2240 61665 2268 61696
rect 2225 61659 2283 61665
rect 2225 61625 2237 61659
rect 2271 61625 2283 61659
rect 2225 61619 2283 61625
rect 1486 61588 1492 61600
rect 1447 61560 1492 61588
rect 1486 61548 1492 61560
rect 1544 61548 1550 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5845 61498
rect 5897 61446 5909 61498
rect 5961 61446 5973 61498
rect 6025 61446 6037 61498
rect 6089 61446 6101 61498
rect 6153 61446 9109 61498
rect 9161 61446 9173 61498
rect 9225 61446 9237 61498
rect 9289 61446 9301 61498
rect 9353 61446 9365 61498
rect 9417 61446 10856 61498
rect 1104 61424 10856 61446
rect 4062 61384 4068 61396
rect 1688 61356 4068 61384
rect 1688 61189 1716 61356
rect 4062 61344 4068 61356
rect 4120 61344 4126 61396
rect 2958 61316 2964 61328
rect 2424 61288 2964 61316
rect 2424 61189 2452 61288
rect 2958 61276 2964 61288
rect 3016 61316 3022 61328
rect 3602 61316 3608 61328
rect 3016 61288 3608 61316
rect 3016 61276 3022 61288
rect 3602 61276 3608 61288
rect 3660 61276 3666 61328
rect 3786 61248 3792 61260
rect 2608 61220 3792 61248
rect 2608 61189 2636 61220
rect 3786 61208 3792 61220
rect 3844 61208 3850 61260
rect 1673 61183 1731 61189
rect 1673 61149 1685 61183
rect 1719 61149 1731 61183
rect 1673 61143 1731 61149
rect 2409 61183 2467 61189
rect 2409 61149 2421 61183
rect 2455 61149 2467 61183
rect 2409 61143 2467 61149
rect 2593 61183 2651 61189
rect 2593 61149 2605 61183
rect 2639 61149 2651 61183
rect 2593 61143 2651 61149
rect 2777 61183 2835 61189
rect 2777 61149 2789 61183
rect 2823 61180 2835 61183
rect 3326 61180 3332 61192
rect 2823 61152 3332 61180
rect 2823 61149 2835 61152
rect 2777 61143 2835 61149
rect 3326 61140 3332 61152
rect 3384 61180 3390 61192
rect 3878 61180 3884 61192
rect 3384 61152 3884 61180
rect 3384 61140 3390 61152
rect 3878 61140 3884 61152
rect 3936 61140 3942 61192
rect 10134 61180 10140 61192
rect 10095 61152 10140 61180
rect 10134 61140 10140 61152
rect 10192 61140 10198 61192
rect 2685 61115 2743 61121
rect 2685 61081 2697 61115
rect 2731 61112 2743 61115
rect 11609 61115 11667 61121
rect 11609 61112 11621 61115
rect 2731 61084 11621 61112
rect 2731 61081 2743 61084
rect 2685 61075 2743 61081
rect 11609 61081 11621 61084
rect 11655 61081 11667 61115
rect 11609 61075 11667 61081
rect 1394 61004 1400 61056
rect 1452 61044 1458 61056
rect 1489 61047 1547 61053
rect 1489 61044 1501 61047
rect 1452 61016 1501 61044
rect 1452 61004 1458 61016
rect 1489 61013 1501 61016
rect 1535 61013 1547 61047
rect 1489 61007 1547 61013
rect 2961 61047 3019 61053
rect 2961 61013 2973 61047
rect 3007 61044 3019 61047
rect 3142 61044 3148 61056
rect 3007 61016 3148 61044
rect 3007 61013 3019 61016
rect 2961 61007 3019 61013
rect 3142 61004 3148 61016
rect 3200 61004 3206 61056
rect 9950 61044 9956 61056
rect 9911 61016 9956 61044
rect 9950 61004 9956 61016
rect 10008 61004 10014 61056
rect 1104 60954 10856 60976
rect 1104 60902 4213 60954
rect 4265 60902 4277 60954
rect 4329 60902 4341 60954
rect 4393 60902 4405 60954
rect 4457 60902 4469 60954
rect 4521 60902 7477 60954
rect 7529 60902 7541 60954
rect 7593 60902 7605 60954
rect 7657 60902 7669 60954
rect 7721 60902 7733 60954
rect 7785 60902 10856 60954
rect 1104 60880 10856 60902
rect 2130 60840 2136 60852
rect 1924 60812 2136 60840
rect 1670 60732 1676 60784
rect 1728 60772 1734 60784
rect 1728 60744 1773 60772
rect 1728 60732 1734 60744
rect 1924 60713 1952 60812
rect 2130 60800 2136 60812
rect 2188 60840 2194 60852
rect 2590 60840 2596 60852
rect 2188 60812 2596 60840
rect 2188 60800 2194 60812
rect 2590 60800 2596 60812
rect 2648 60800 2654 60852
rect 9858 60772 9864 60784
rect 2700 60744 9864 60772
rect 1535 60707 1593 60713
rect 1535 60673 1547 60707
rect 1581 60704 1593 60707
rect 1765 60707 1823 60713
rect 1581 60676 1716 60704
rect 1581 60673 1593 60676
rect 1535 60667 1593 60673
rect 1688 60648 1716 60676
rect 1765 60673 1777 60707
rect 1811 60673 1823 60707
rect 1765 60667 1823 60673
rect 1909 60707 1967 60713
rect 1909 60673 1921 60707
rect 1955 60673 1967 60707
rect 2593 60707 2651 60713
rect 2593 60704 2605 60707
rect 1909 60667 1967 60673
rect 2240 60676 2605 60704
rect 1670 60596 1676 60648
rect 1728 60596 1734 60648
rect 1780 60568 1808 60667
rect 2240 60648 2268 60676
rect 2593 60673 2605 60676
rect 2639 60673 2651 60707
rect 2593 60667 2651 60673
rect 2222 60596 2228 60648
rect 2280 60596 2286 60648
rect 2700 60568 2728 60744
rect 9858 60732 9864 60744
rect 9916 60732 9922 60784
rect 10134 60704 10140 60716
rect 10095 60676 10140 60704
rect 10134 60664 10140 60676
rect 10192 60664 10198 60716
rect 1780 60540 2728 60568
rect 2774 60528 2780 60580
rect 2832 60568 2838 60580
rect 2832 60540 2877 60568
rect 2832 60528 2838 60540
rect 474 60460 480 60512
rect 532 60500 538 60512
rect 1210 60500 1216 60512
rect 532 60472 1216 60500
rect 532 60460 538 60472
rect 1210 60460 1216 60472
rect 1268 60460 1274 60512
rect 2041 60503 2099 60509
rect 2041 60469 2053 60503
rect 2087 60500 2099 60503
rect 6362 60500 6368 60512
rect 2087 60472 6368 60500
rect 2087 60469 2099 60472
rect 2041 60463 2099 60469
rect 6362 60460 6368 60472
rect 6420 60460 6426 60512
rect 9950 60500 9956 60512
rect 9911 60472 9956 60500
rect 9950 60460 9956 60472
rect 10008 60460 10014 60512
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5845 60410
rect 5897 60358 5909 60410
rect 5961 60358 5973 60410
rect 6025 60358 6037 60410
rect 6089 60358 6101 60410
rect 6153 60358 9109 60410
rect 9161 60358 9173 60410
rect 9225 60358 9237 60410
rect 9289 60358 9301 60410
rect 9353 60358 9365 60410
rect 9417 60358 10856 60410
rect 1104 60336 10856 60358
rect 2498 60256 2504 60308
rect 2556 60296 2562 60308
rect 2556 60268 2774 60296
rect 2556 60256 2562 60268
rect 1210 60188 1216 60240
rect 1268 60228 1274 60240
rect 2593 60231 2651 60237
rect 2593 60228 2605 60231
rect 1268 60200 2605 60228
rect 1268 60188 1274 60200
rect 2593 60197 2605 60200
rect 2639 60197 2651 60231
rect 2593 60191 2651 60197
rect 845 60095 903 60101
rect 845 60061 857 60095
rect 891 60092 903 60095
rect 1670 60092 1676 60104
rect 891 60064 1676 60092
rect 891 60061 903 60064
rect 845 60055 903 60061
rect 1670 60052 1676 60064
rect 1728 60092 1734 60104
rect 2041 60095 2099 60101
rect 2041 60092 2053 60095
rect 1728 60064 2053 60092
rect 1728 60052 1734 60064
rect 2041 60061 2053 60064
rect 2087 60061 2099 60095
rect 2041 60055 2099 60061
rect 2461 60095 2519 60101
rect 2461 60061 2473 60095
rect 2507 60092 2519 60095
rect 2590 60092 2596 60104
rect 2507 60064 2596 60092
rect 2507 60061 2519 60064
rect 2461 60055 2519 60061
rect 2590 60052 2596 60064
rect 2648 60092 2654 60104
rect 2746 60092 2774 60268
rect 2648 60064 2774 60092
rect 2648 60052 2654 60064
rect 2225 60027 2283 60033
rect 2225 59993 2237 60027
rect 2271 59993 2283 60027
rect 2225 59987 2283 59993
rect 2317 60027 2375 60033
rect 2317 59993 2329 60027
rect 2363 60024 2375 60027
rect 9858 60024 9864 60036
rect 2363 59996 9864 60024
rect 2363 59993 2375 59996
rect 2317 59987 2375 59993
rect 2240 59956 2268 59987
rect 9858 59984 9864 59996
rect 9916 59984 9922 60036
rect 3510 59956 3516 59968
rect 2240 59928 3516 59956
rect 3510 59916 3516 59928
rect 3568 59916 3574 59968
rect 1104 59866 10856 59888
rect 1104 59814 4213 59866
rect 4265 59814 4277 59866
rect 4329 59814 4341 59866
rect 4393 59814 4405 59866
rect 4457 59814 4469 59866
rect 4521 59814 7477 59866
rect 7529 59814 7541 59866
rect 7593 59814 7605 59866
rect 7657 59814 7669 59866
rect 7721 59814 7733 59866
rect 7785 59814 10856 59866
rect 1104 59792 10856 59814
rect 1670 59712 1676 59764
rect 1728 59712 1734 59764
rect 1688 59684 1716 59712
rect 2314 59684 2320 59696
rect 1688 59656 2176 59684
rect 2275 59656 2320 59684
rect 2148 59625 2176 59656
rect 2314 59644 2320 59656
rect 2372 59644 2378 59696
rect 2409 59687 2467 59693
rect 2409 59653 2421 59687
rect 2455 59684 2467 59687
rect 9766 59684 9772 59696
rect 2455 59656 9772 59684
rect 2455 59653 2467 59656
rect 2409 59647 2467 59653
rect 9766 59644 9772 59656
rect 9824 59644 9830 59696
rect 2590 59625 2596 59628
rect 1673 59619 1731 59625
rect 1673 59585 1685 59619
rect 1719 59585 1731 59619
rect 1673 59579 1731 59585
rect 2133 59619 2191 59625
rect 2133 59585 2145 59619
rect 2179 59585 2191 59619
rect 2553 59619 2596 59625
rect 2553 59616 2565 59619
rect 2133 59579 2191 59585
rect 2332 59588 2565 59616
rect 1688 59480 1716 59579
rect 2332 59560 2360 59588
rect 2553 59585 2565 59588
rect 2553 59579 2596 59585
rect 2590 59576 2596 59579
rect 2648 59576 2654 59628
rect 2682 59576 2688 59628
rect 2740 59616 2746 59628
rect 3237 59619 3295 59625
rect 3237 59616 3249 59619
rect 2740 59588 3249 59616
rect 2740 59576 2746 59588
rect 3237 59585 3249 59588
rect 3283 59585 3295 59619
rect 10134 59616 10140 59628
rect 10095 59588 10140 59616
rect 3237 59579 3295 59585
rect 10134 59576 10140 59588
rect 10192 59576 10198 59628
rect 2314 59508 2320 59560
rect 2372 59508 2378 59560
rect 4982 59548 4988 59560
rect 2746 59520 4988 59548
rect 2746 59480 2774 59520
rect 4982 59508 4988 59520
rect 5040 59508 5046 59560
rect 1688 59452 2774 59480
rect 3050 59440 3056 59492
rect 3108 59480 3114 59492
rect 3421 59483 3479 59489
rect 3421 59480 3433 59483
rect 3108 59452 3433 59480
rect 3108 59440 3114 59452
rect 3421 59449 3433 59452
rect 3467 59449 3479 59483
rect 3421 59443 3479 59449
rect 1486 59412 1492 59424
rect 1447 59384 1492 59412
rect 1486 59372 1492 59384
rect 1544 59372 1550 59424
rect 2685 59415 2743 59421
rect 2685 59381 2697 59415
rect 2731 59412 2743 59415
rect 3234 59412 3240 59424
rect 2731 59384 3240 59412
rect 2731 59381 2743 59384
rect 2685 59375 2743 59381
rect 3234 59372 3240 59384
rect 3292 59372 3298 59424
rect 9953 59415 10011 59421
rect 9953 59381 9965 59415
rect 9999 59412 10011 59415
rect 11517 59415 11575 59421
rect 11517 59412 11529 59415
rect 9999 59384 11529 59412
rect 9999 59381 10011 59384
rect 9953 59375 10011 59381
rect 11517 59381 11529 59384
rect 11563 59381 11575 59415
rect 11517 59375 11575 59381
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5845 59322
rect 5897 59270 5909 59322
rect 5961 59270 5973 59322
rect 6025 59270 6037 59322
rect 6089 59270 6101 59322
rect 6153 59270 9109 59322
rect 9161 59270 9173 59322
rect 9225 59270 9237 59322
rect 9289 59270 9301 59322
rect 9353 59270 9365 59322
rect 9417 59270 10856 59322
rect 1104 59248 10856 59270
rect 1394 59168 1400 59220
rect 1452 59208 1458 59220
rect 2593 59211 2651 59217
rect 2593 59208 2605 59211
rect 1452 59180 2605 59208
rect 1452 59168 1458 59180
rect 2593 59177 2605 59180
rect 2639 59177 2651 59211
rect 2593 59171 2651 59177
rect 753 59143 811 59149
rect 753 59109 765 59143
rect 799 59140 811 59143
rect 1578 59140 1584 59152
rect 799 59112 1584 59140
rect 799 59109 811 59112
rect 753 59103 811 59109
rect 1578 59100 1584 59112
rect 1636 59100 1642 59152
rect 1949 59143 2007 59149
rect 1949 59109 1961 59143
rect 1995 59140 2007 59143
rect 11885 59143 11943 59149
rect 11885 59140 11897 59143
rect 1995 59112 11897 59140
rect 1995 59109 2007 59112
rect 1949 59103 2007 59109
rect 11885 59109 11897 59112
rect 11931 59109 11943 59143
rect 11885 59103 11943 59109
rect 1670 59072 1676 59084
rect 1412 59044 1676 59072
rect 1412 59013 1440 59044
rect 1670 59032 1676 59044
rect 1728 59032 1734 59084
rect 1397 59007 1455 59013
rect 1397 58973 1409 59007
rect 1443 58973 1455 59007
rect 1578 59004 1584 59016
rect 1539 58976 1584 59004
rect 1397 58967 1455 58973
rect 1302 58828 1308 58880
rect 1360 58868 1366 58880
rect 1412 58868 1440 58967
rect 1578 58964 1584 58976
rect 1636 58964 1642 59016
rect 1817 59007 1875 59013
rect 1817 58973 1829 59007
rect 1863 59004 1875 59007
rect 2314 59004 2320 59016
rect 1863 58976 2320 59004
rect 1863 58973 1875 58976
rect 1817 58967 1875 58973
rect 2314 58964 2320 58976
rect 2372 58964 2378 59016
rect 2777 59007 2835 59013
rect 2777 58973 2789 59007
rect 2823 59004 2835 59007
rect 3786 59004 3792 59016
rect 2823 58976 3792 59004
rect 2823 58973 2835 58976
rect 2777 58967 2835 58973
rect 3786 58964 3792 58976
rect 3844 58964 3850 59016
rect 9950 58964 9956 59016
rect 10008 58964 10014 59016
rect 10134 59004 10140 59016
rect 10095 58976 10140 59004
rect 10134 58964 10140 58976
rect 10192 58964 10198 59016
rect 1673 58939 1731 58945
rect 1673 58905 1685 58939
rect 1719 58936 1731 58939
rect 9968 58936 9996 58964
rect 1719 58908 9996 58936
rect 1719 58905 1731 58908
rect 1673 58899 1731 58905
rect 9950 58868 9956 58880
rect 1360 58840 1440 58868
rect 9911 58840 9956 58868
rect 1360 58828 1366 58840
rect 9950 58828 9956 58840
rect 10008 58828 10014 58880
rect 1104 58778 10856 58800
rect 1104 58726 4213 58778
rect 4265 58726 4277 58778
rect 4329 58726 4341 58778
rect 4393 58726 4405 58778
rect 4457 58726 4469 58778
rect 4521 58726 7477 58778
rect 7529 58726 7541 58778
rect 7593 58726 7605 58778
rect 7657 58726 7669 58778
rect 7721 58726 7733 58778
rect 7785 58726 10856 58778
rect 1104 58704 10856 58726
rect 658 58624 664 58676
rect 716 58664 722 58676
rect 716 58636 2636 58664
rect 716 58624 722 58636
rect 1857 58599 1915 58605
rect 1857 58565 1869 58599
rect 1903 58596 1915 58599
rect 1903 58568 2360 58596
rect 1903 58565 1915 58568
rect 1857 58559 1915 58565
rect 1670 58488 1676 58540
rect 1728 58537 1734 58540
rect 1728 58531 1771 58537
rect 1759 58497 1771 58531
rect 1946 58528 1952 58540
rect 1907 58500 1952 58528
rect 1728 58491 1771 58497
rect 1728 58488 1734 58491
rect 1946 58488 1952 58500
rect 2004 58488 2010 58540
rect 2133 58531 2191 58537
rect 2133 58497 2145 58531
rect 2179 58497 2191 58531
rect 2133 58491 2191 58497
rect 1302 58420 1308 58472
rect 1360 58460 1366 58472
rect 2148 58460 2176 58491
rect 1360 58432 2176 58460
rect 2332 58460 2360 58568
rect 2608 58537 2636 58636
rect 11057 58599 11115 58605
rect 11057 58596 11069 58599
rect 2746 58568 11069 58596
rect 2593 58531 2651 58537
rect 2593 58497 2605 58531
rect 2639 58497 2651 58531
rect 2593 58491 2651 58497
rect 2746 58460 2774 58568
rect 11057 58565 11069 58568
rect 11103 58565 11115 58599
rect 11057 58559 11115 58565
rect 9861 58531 9919 58537
rect 9861 58497 9873 58531
rect 9907 58528 9919 58531
rect 11793 58531 11851 58537
rect 11793 58528 11805 58531
rect 9907 58500 11805 58528
rect 9907 58497 9919 58500
rect 9861 58491 9919 58497
rect 11793 58497 11805 58500
rect 11839 58497 11851 58531
rect 11793 58491 11851 58497
rect 10134 58460 10140 58472
rect 2332 58432 2774 58460
rect 10095 58432 10140 58460
rect 1360 58420 1366 58432
rect 10134 58420 10140 58432
rect 10192 58420 10198 58472
rect 8570 58392 8576 58404
rect 2148 58364 8576 58392
rect 1581 58327 1639 58333
rect 1581 58293 1593 58327
rect 1627 58324 1639 58327
rect 2148 58324 2176 58364
rect 8570 58352 8576 58364
rect 8628 58352 8634 58404
rect 1627 58296 2176 58324
rect 1627 58293 1639 58296
rect 1581 58287 1639 58293
rect 2406 58284 2412 58336
rect 2464 58324 2470 58336
rect 2777 58327 2835 58333
rect 2777 58324 2789 58327
rect 2464 58296 2789 58324
rect 2464 58284 2470 58296
rect 2777 58293 2789 58296
rect 2823 58293 2835 58327
rect 2777 58287 2835 58293
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5845 58234
rect 5897 58182 5909 58234
rect 5961 58182 5973 58234
rect 6025 58182 6037 58234
rect 6089 58182 6101 58234
rect 6153 58182 9109 58234
rect 9161 58182 9173 58234
rect 9225 58182 9237 58234
rect 9289 58182 9301 58234
rect 9353 58182 9365 58234
rect 9417 58182 10856 58234
rect 1104 58160 10856 58182
rect 2406 58052 2412 58064
rect 1596 58024 2412 58052
rect 1302 57944 1308 57996
rect 1360 57984 1366 57996
rect 1596 57984 1624 58024
rect 2406 58012 2412 58024
rect 2464 58012 2470 58064
rect 3510 58012 3516 58064
rect 3568 58052 3574 58064
rect 4062 58052 4068 58064
rect 3568 58024 4068 58052
rect 3568 58012 3574 58024
rect 4062 58012 4068 58024
rect 4120 58012 4126 58064
rect 1360 57956 1624 57984
rect 1360 57944 1366 57956
rect 1489 57919 1547 57925
rect 1489 57885 1501 57919
rect 1535 57916 1547 57919
rect 1596 57916 1624 57956
rect 1670 57944 1676 57996
rect 1728 57944 1734 57996
rect 2516 57956 2774 57984
rect 1535 57888 1624 57916
rect 1688 57916 1716 57944
rect 1946 57925 1952 57928
rect 1909 57919 1952 57925
rect 1909 57916 1921 57919
rect 1688 57888 1921 57916
rect 1535 57885 1547 57888
rect 1489 57879 1547 57885
rect 1909 57885 1921 57888
rect 1909 57879 1952 57885
rect 1946 57876 1952 57879
rect 2004 57876 2010 57928
rect 2058 57919 2116 57925
rect 2058 57885 2070 57919
rect 2104 57916 2116 57919
rect 2516 57916 2544 57956
rect 2104 57888 2544 57916
rect 2104 57885 2116 57888
rect 2058 57879 2116 57885
rect 2590 57876 2596 57928
rect 2648 57916 2654 57928
rect 2746 57916 2774 57956
rect 3050 57916 3056 57928
rect 2648 57888 2693 57916
rect 2746 57888 3056 57916
rect 2648 57876 2654 57888
rect 3050 57876 3056 57888
rect 3108 57876 3114 57928
rect 3878 57916 3884 57928
rect 3839 57888 3884 57916
rect 3878 57876 3884 57888
rect 3936 57876 3942 57928
rect 3973 57919 4031 57925
rect 3973 57885 3985 57919
rect 4019 57916 4031 57919
rect 4062 57916 4068 57928
rect 4019 57888 4068 57916
rect 4019 57885 4031 57888
rect 3973 57879 4031 57885
rect 4062 57876 4068 57888
rect 4120 57876 4126 57928
rect 1673 57851 1731 57857
rect 1673 57817 1685 57851
rect 1719 57817 1731 57851
rect 1673 57811 1731 57817
rect 1765 57851 1823 57857
rect 1765 57817 1777 57851
rect 1811 57848 1823 57851
rect 9950 57848 9956 57860
rect 1811 57820 9956 57848
rect 1811 57817 1823 57820
rect 1765 57811 1823 57817
rect 1688 57780 1716 57811
rect 9950 57808 9956 57820
rect 10008 57808 10014 57860
rect 2314 57780 2320 57792
rect 1688 57752 2320 57780
rect 2314 57740 2320 57752
rect 2372 57740 2378 57792
rect 2774 57740 2780 57792
rect 2832 57780 2838 57792
rect 2832 57752 2877 57780
rect 2832 57740 2838 57752
rect 3234 57740 3240 57792
rect 3292 57780 3298 57792
rect 3878 57780 3884 57792
rect 3292 57752 3884 57780
rect 3292 57740 3298 57752
rect 3878 57740 3884 57752
rect 3936 57740 3942 57792
rect 1104 57690 10856 57712
rect 1104 57638 4213 57690
rect 4265 57638 4277 57690
rect 4329 57638 4341 57690
rect 4393 57638 4405 57690
rect 4457 57638 4469 57690
rect 4521 57638 7477 57690
rect 7529 57638 7541 57690
rect 7593 57638 7605 57690
rect 7657 57638 7669 57690
rect 7721 57638 7733 57690
rect 7785 57638 10856 57690
rect 1104 57616 10856 57638
rect 106 57536 112 57588
rect 164 57576 170 57588
rect 2590 57576 2596 57588
rect 164 57548 2596 57576
rect 164 57536 170 57548
rect 2590 57536 2596 57548
rect 2648 57536 2654 57588
rect 2961 57579 3019 57585
rect 2961 57545 2973 57579
rect 3007 57576 3019 57579
rect 3326 57576 3332 57588
rect 3007 57548 3332 57576
rect 3007 57545 3019 57548
rect 2961 57539 3019 57545
rect 3326 57536 3332 57548
rect 3384 57536 3390 57588
rect 4890 57508 4896 57520
rect 2746 57480 4896 57508
rect 1673 57443 1731 57449
rect 1673 57409 1685 57443
rect 1719 57409 1731 57443
rect 1673 57403 1731 57409
rect 2409 57443 2467 57449
rect 2409 57409 2421 57443
rect 2455 57440 2467 57443
rect 2746 57440 2774 57480
rect 4890 57468 4896 57480
rect 4948 57468 4954 57520
rect 2455 57412 2774 57440
rect 2869 57443 2927 57449
rect 2455 57409 2467 57412
rect 2409 57403 2467 57409
rect 2869 57409 2881 57443
rect 2915 57409 2927 57443
rect 2869 57403 2927 57409
rect 3053 57443 3111 57449
rect 3053 57409 3065 57443
rect 3099 57440 3111 57443
rect 3234 57440 3240 57452
rect 3099 57412 3240 57440
rect 3099 57409 3111 57412
rect 3053 57403 3111 57409
rect 1486 57236 1492 57248
rect 1447 57208 1492 57236
rect 1486 57196 1492 57208
rect 1544 57196 1550 57248
rect 1688 57236 1716 57403
rect 2884 57372 2912 57403
rect 3234 57400 3240 57412
rect 3292 57400 3298 57452
rect 9861 57443 9919 57449
rect 9861 57409 9873 57443
rect 9907 57440 9919 57443
rect 11609 57443 11667 57449
rect 11609 57440 11621 57443
rect 9907 57412 11621 57440
rect 9907 57409 9919 57412
rect 9861 57403 9919 57409
rect 11609 57409 11621 57412
rect 11655 57409 11667 57443
rect 11609 57403 11667 57409
rect 3326 57372 3332 57384
rect 2884 57344 3332 57372
rect 3326 57332 3332 57344
rect 3384 57332 3390 57384
rect 10134 57372 10140 57384
rect 10095 57344 10140 57372
rect 10134 57332 10140 57344
rect 10192 57332 10198 57384
rect 2222 57304 2228 57316
rect 2183 57276 2228 57304
rect 2222 57264 2228 57276
rect 2280 57264 2286 57316
rect 5350 57236 5356 57248
rect 1688 57208 5356 57236
rect 5350 57196 5356 57208
rect 5408 57196 5414 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5845 57146
rect 5897 57094 5909 57146
rect 5961 57094 5973 57146
rect 6025 57094 6037 57146
rect 6089 57094 6101 57146
rect 6153 57094 9109 57146
rect 9161 57094 9173 57146
rect 9225 57094 9237 57146
rect 9289 57094 9301 57146
rect 9353 57094 9365 57146
rect 9417 57094 10856 57146
rect 1104 57072 10856 57094
rect 2958 56992 2964 57044
rect 3016 57032 3022 57044
rect 3053 57035 3111 57041
rect 3053 57032 3065 57035
rect 3016 57004 3065 57032
rect 3016 56992 3022 57004
rect 3053 57001 3065 57004
rect 3099 57001 3111 57035
rect 3053 56995 3111 57001
rect 2406 56924 2412 56976
rect 2464 56964 2470 56976
rect 2590 56964 2596 56976
rect 2464 56936 2596 56964
rect 2464 56924 2470 56936
rect 2590 56924 2596 56936
rect 2648 56924 2654 56976
rect 6638 56896 6644 56908
rect 3804 56868 6644 56896
rect 750 56788 756 56840
rect 808 56828 814 56840
rect 1673 56831 1731 56837
rect 1673 56828 1685 56831
rect 808 56800 1685 56828
rect 808 56788 814 56800
rect 1673 56797 1685 56800
rect 1719 56797 1731 56831
rect 2406 56828 2412 56840
rect 2367 56800 2412 56828
rect 1673 56791 1731 56797
rect 2406 56788 2412 56800
rect 2464 56788 2470 56840
rect 2869 56831 2927 56837
rect 2869 56797 2881 56831
rect 2915 56797 2927 56831
rect 2869 56791 2927 56797
rect 3053 56831 3111 56837
rect 3053 56797 3065 56831
rect 3099 56828 3111 56831
rect 3326 56828 3332 56840
rect 3099 56800 3332 56828
rect 3099 56797 3111 56800
rect 3053 56791 3111 56797
rect 2884 56760 2912 56791
rect 3326 56788 3332 56800
rect 3384 56788 3390 56840
rect 3804 56837 3832 56868
rect 6638 56856 6644 56868
rect 6696 56856 6702 56908
rect 9861 56899 9919 56905
rect 9861 56865 9873 56899
rect 9907 56896 9919 56899
rect 11701 56899 11759 56905
rect 11701 56896 11713 56899
rect 9907 56868 11713 56896
rect 9907 56865 9919 56868
rect 9861 56859 9919 56865
rect 11701 56865 11713 56868
rect 11747 56865 11759 56899
rect 11701 56859 11759 56865
rect 3789 56831 3847 56837
rect 3789 56828 3801 56831
rect 3436 56800 3801 56828
rect 3436 56760 3464 56800
rect 3789 56797 3801 56800
rect 3835 56797 3847 56831
rect 3789 56791 3847 56797
rect 3973 56831 4031 56837
rect 3973 56797 3985 56831
rect 4019 56828 4031 56831
rect 4062 56828 4068 56840
rect 4019 56800 4068 56828
rect 4019 56797 4031 56800
rect 3973 56791 4031 56797
rect 2884 56732 3464 56760
rect 3510 56720 3516 56772
rect 3568 56760 3574 56772
rect 3988 56760 4016 56791
rect 4062 56788 4068 56800
rect 4120 56788 4126 56840
rect 10134 56828 10140 56840
rect 10095 56800 10140 56828
rect 10134 56788 10140 56800
rect 10192 56788 10198 56840
rect 3568 56732 4016 56760
rect 3568 56720 3574 56732
rect 1486 56692 1492 56704
rect 1447 56664 1492 56692
rect 1486 56652 1492 56664
rect 1544 56652 1550 56704
rect 2222 56692 2228 56704
rect 2183 56664 2228 56692
rect 2222 56652 2228 56664
rect 2280 56652 2286 56704
rect 3881 56695 3939 56701
rect 3881 56661 3893 56695
rect 3927 56692 3939 56695
rect 11057 56695 11115 56701
rect 11057 56692 11069 56695
rect 3927 56664 11069 56692
rect 3927 56661 3939 56664
rect 3881 56655 3939 56661
rect 11057 56661 11069 56664
rect 11103 56661 11115 56695
rect 11057 56655 11115 56661
rect 1104 56602 10856 56624
rect 1104 56550 4213 56602
rect 4265 56550 4277 56602
rect 4329 56550 4341 56602
rect 4393 56550 4405 56602
rect 4457 56550 4469 56602
rect 4521 56550 7477 56602
rect 7529 56550 7541 56602
rect 7593 56550 7605 56602
rect 7657 56550 7669 56602
rect 7721 56550 7733 56602
rect 7785 56550 10856 56602
rect 1104 56528 10856 56550
rect 1394 56448 1400 56500
rect 1452 56488 1458 56500
rect 1670 56488 1676 56500
rect 1452 56460 1676 56488
rect 1452 56448 1458 56460
rect 1670 56448 1676 56460
rect 1728 56448 1734 56500
rect 8846 56488 8852 56500
rect 2746 56460 8852 56488
rect 753 56423 811 56429
rect 753 56389 765 56423
rect 799 56420 811 56423
rect 2590 56420 2596 56432
rect 799 56392 2596 56420
rect 799 56389 811 56392
rect 753 56383 811 56389
rect 2590 56380 2596 56392
rect 2648 56380 2654 56432
rect 1673 56355 1731 56361
rect 1673 56321 1685 56355
rect 1719 56352 1731 56355
rect 2746 56352 2774 56460
rect 8846 56448 8852 56460
rect 8904 56448 8910 56500
rect 2958 56420 2964 56432
rect 2871 56392 2964 56420
rect 2884 56361 2912 56392
rect 2958 56380 2964 56392
rect 3016 56420 3022 56432
rect 3602 56420 3608 56432
rect 3016 56392 3608 56420
rect 3016 56380 3022 56392
rect 3602 56380 3608 56392
rect 3660 56380 3666 56432
rect 1719 56324 2774 56352
rect 2869 56355 2927 56361
rect 1719 56321 1731 56324
rect 1673 56315 1731 56321
rect 2869 56321 2881 56355
rect 2915 56321 2927 56355
rect 2869 56315 2927 56321
rect 3234 56312 3240 56364
rect 3292 56352 3298 56364
rect 3329 56355 3387 56361
rect 3329 56352 3341 56355
rect 3292 56324 3341 56352
rect 3292 56312 3298 56324
rect 3329 56321 3341 56324
rect 3375 56321 3387 56355
rect 3510 56352 3516 56364
rect 3471 56324 3516 56352
rect 3329 56315 3387 56321
rect 1394 56244 1400 56296
rect 1452 56284 1458 56296
rect 1946 56284 1952 56296
rect 1452 56256 1952 56284
rect 1452 56244 1458 56256
rect 1946 56244 1952 56256
rect 2004 56244 2010 56296
rect 3344 56284 3372 56315
rect 3510 56312 3516 56324
rect 3568 56312 3574 56364
rect 5258 56284 5264 56296
rect 3344 56256 5264 56284
rect 5258 56244 5264 56256
rect 5316 56244 5322 56296
rect 3234 56176 3240 56228
rect 3292 56216 3298 56228
rect 3878 56216 3884 56228
rect 3292 56188 3884 56216
rect 3292 56176 3298 56188
rect 3878 56176 3884 56188
rect 3936 56176 3942 56228
rect 1394 56108 1400 56160
rect 1452 56148 1458 56160
rect 1489 56151 1547 56157
rect 1489 56148 1501 56151
rect 1452 56120 1501 56148
rect 1452 56108 1458 56120
rect 1489 56117 1501 56120
rect 1535 56117 1547 56151
rect 1489 56111 1547 56117
rect 1946 56108 1952 56160
rect 2004 56148 2010 56160
rect 2130 56148 2136 56160
rect 2004 56120 2136 56148
rect 2004 56108 2010 56120
rect 2130 56108 2136 56120
rect 2188 56108 2194 56160
rect 3513 56151 3571 56157
rect 3513 56117 3525 56151
rect 3559 56148 3571 56151
rect 9858 56148 9864 56160
rect 3559 56120 9864 56148
rect 3559 56117 3571 56120
rect 3513 56111 3571 56117
rect 9858 56108 9864 56120
rect 9916 56108 9922 56160
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5845 56058
rect 5897 56006 5909 56058
rect 5961 56006 5973 56058
rect 6025 56006 6037 56058
rect 6089 56006 6101 56058
rect 6153 56006 9109 56058
rect 9161 56006 9173 56058
rect 9225 56006 9237 56058
rect 9289 56006 9301 56058
rect 9353 56006 9365 56058
rect 9417 56006 10856 56058
rect 1104 55984 10856 56006
rect 2958 55944 2964 55956
rect 2919 55916 2964 55944
rect 2958 55904 2964 55916
rect 3016 55904 3022 55956
rect 4798 55876 4804 55888
rect 1688 55848 4804 55876
rect 1688 55749 1716 55848
rect 4798 55836 4804 55848
rect 4856 55836 4862 55888
rect 8754 55808 8760 55820
rect 2148 55780 8760 55808
rect 2148 55749 2176 55780
rect 8754 55768 8760 55780
rect 8812 55768 8818 55820
rect 1673 55743 1731 55749
rect 1673 55709 1685 55743
rect 1719 55709 1731 55743
rect 1673 55703 1731 55709
rect 2133 55743 2191 55749
rect 2133 55709 2145 55743
rect 2179 55709 2191 55743
rect 3050 55740 3056 55752
rect 3011 55712 3056 55740
rect 2133 55703 2191 55709
rect 3050 55700 3056 55712
rect 3108 55700 3114 55752
rect 10134 55740 10140 55752
rect 10095 55712 10140 55740
rect 10134 55700 10140 55712
rect 10192 55700 10198 55752
rect 1486 55604 1492 55616
rect 1447 55576 1492 55604
rect 1486 55564 1492 55576
rect 1544 55564 1550 55616
rect 2314 55604 2320 55616
rect 2275 55576 2320 55604
rect 2314 55564 2320 55576
rect 2372 55564 2378 55616
rect 9953 55607 10011 55613
rect 9953 55573 9965 55607
rect 9999 55604 10011 55607
rect 11241 55607 11299 55613
rect 11241 55604 11253 55607
rect 9999 55576 11253 55604
rect 9999 55573 10011 55576
rect 9953 55567 10011 55573
rect 11241 55573 11253 55576
rect 11287 55573 11299 55607
rect 11241 55567 11299 55573
rect 1104 55514 10856 55536
rect 1104 55462 4213 55514
rect 4265 55462 4277 55514
rect 4329 55462 4341 55514
rect 4393 55462 4405 55514
rect 4457 55462 4469 55514
rect 4521 55462 7477 55514
rect 7529 55462 7541 55514
rect 7593 55462 7605 55514
rect 7657 55462 7669 55514
rect 7721 55462 7733 55514
rect 7785 55462 10856 55514
rect 1104 55440 10856 55462
rect 937 55403 995 55409
rect 937 55369 949 55403
rect 983 55400 995 55403
rect 1210 55400 1216 55412
rect 983 55372 1216 55400
rect 983 55369 995 55372
rect 937 55363 995 55369
rect 1210 55360 1216 55372
rect 1268 55360 1274 55412
rect 11517 55403 11575 55409
rect 11517 55400 11529 55403
rect 1688 55372 11529 55400
rect 1578 55332 1584 55344
rect 1539 55304 1584 55332
rect 1578 55292 1584 55304
rect 1636 55292 1642 55344
rect 1688 55341 1716 55372
rect 11517 55369 11529 55372
rect 11563 55369 11575 55403
rect 11517 55363 11575 55369
rect 1673 55335 1731 55341
rect 1673 55301 1685 55335
rect 1719 55301 1731 55335
rect 3326 55332 3332 55344
rect 3287 55304 3332 55332
rect 1673 55295 1731 55301
rect 3326 55292 3332 55304
rect 3384 55292 3390 55344
rect 753 55267 811 55273
rect 753 55233 765 55267
rect 799 55264 811 55267
rect 1397 55267 1455 55273
rect 1397 55264 1409 55267
rect 799 55236 1409 55264
rect 799 55233 811 55236
rect 753 55227 811 55233
rect 1397 55233 1409 55236
rect 1443 55233 1455 55267
rect 1765 55267 1823 55273
rect 1765 55264 1777 55267
rect 1397 55227 1455 55233
rect 1596 55236 1777 55264
rect 1596 55208 1624 55236
rect 1765 55233 1777 55236
rect 1811 55233 1823 55267
rect 1765 55227 1823 55233
rect 2314 55224 2320 55276
rect 2372 55264 2378 55276
rect 2593 55267 2651 55273
rect 2593 55264 2605 55267
rect 2372 55236 2605 55264
rect 2372 55224 2378 55236
rect 2593 55233 2605 55236
rect 2639 55264 2651 55267
rect 3050 55264 3056 55276
rect 2639 55236 3056 55264
rect 2639 55233 2651 55236
rect 2593 55227 2651 55233
rect 3050 55224 3056 55236
rect 3108 55224 3114 55276
rect 10137 55267 10195 55273
rect 10137 55233 10149 55267
rect 10183 55264 10195 55267
rect 10183 55236 10272 55264
rect 10183 55233 10195 55236
rect 10137 55227 10195 55233
rect 10244 55208 10272 55236
rect 1578 55156 1584 55208
rect 1636 55156 1642 55208
rect 10226 55156 10232 55208
rect 10284 55156 10290 55208
rect 1949 55063 2007 55069
rect 1949 55029 1961 55063
rect 1995 55060 2007 55063
rect 2038 55060 2044 55072
rect 1995 55032 2044 55060
rect 1995 55029 2007 55032
rect 1949 55023 2007 55029
rect 2038 55020 2044 55032
rect 2096 55020 2102 55072
rect 9950 55060 9956 55072
rect 9911 55032 9956 55060
rect 9950 55020 9956 55032
rect 10008 55020 10014 55072
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5845 54970
rect 5897 54918 5909 54970
rect 5961 54918 5973 54970
rect 6025 54918 6037 54970
rect 6089 54918 6101 54970
rect 6153 54918 9109 54970
rect 9161 54918 9173 54970
rect 9225 54918 9237 54970
rect 9289 54918 9301 54970
rect 9353 54918 9365 54970
rect 9417 54918 10856 54970
rect 1104 54896 10856 54918
rect 1210 54816 1216 54868
rect 1268 54856 1274 54868
rect 2314 54856 2320 54868
rect 1268 54828 2320 54856
rect 1268 54816 1274 54828
rect 2314 54816 2320 54828
rect 2372 54816 2378 54868
rect 474 54748 480 54800
rect 532 54788 538 54800
rect 3602 54788 3608 54800
rect 532 54760 3608 54788
rect 532 54748 538 54760
rect 3602 54748 3608 54760
rect 3660 54748 3666 54800
rect 1673 54655 1731 54661
rect 1673 54621 1685 54655
rect 1719 54621 1731 54655
rect 1673 54615 1731 54621
rect 2133 54655 2191 54661
rect 2133 54621 2145 54655
rect 2179 54652 2191 54655
rect 4706 54652 4712 54664
rect 2179 54624 4712 54652
rect 2179 54621 2191 54624
rect 2133 54615 2191 54621
rect 1688 54584 1716 54615
rect 4706 54612 4712 54624
rect 4764 54612 4770 54664
rect 5442 54584 5448 54596
rect 1688 54556 5448 54584
rect 5442 54544 5448 54556
rect 5500 54544 5506 54596
rect 1394 54476 1400 54528
rect 1452 54516 1458 54528
rect 1489 54519 1547 54525
rect 1489 54516 1501 54519
rect 1452 54488 1501 54516
rect 1452 54476 1458 54488
rect 1489 54485 1501 54488
rect 1535 54485 1547 54519
rect 1489 54479 1547 54485
rect 2317 54519 2375 54525
rect 2317 54485 2329 54519
rect 2363 54516 2375 54519
rect 2774 54516 2780 54528
rect 2363 54488 2780 54516
rect 2363 54485 2375 54488
rect 2317 54479 2375 54485
rect 2774 54476 2780 54488
rect 2832 54476 2838 54528
rect 1104 54426 10856 54448
rect 1104 54374 4213 54426
rect 4265 54374 4277 54426
rect 4329 54374 4341 54426
rect 4393 54374 4405 54426
rect 4457 54374 4469 54426
rect 4521 54374 7477 54426
rect 7529 54374 7541 54426
rect 7593 54374 7605 54426
rect 7657 54374 7669 54426
rect 7721 54374 7733 54426
rect 7785 54374 10856 54426
rect 1104 54352 10856 54374
rect 1673 54179 1731 54185
rect 1673 54145 1685 54179
rect 1719 54145 1731 54179
rect 1673 54139 1731 54145
rect 2777 54179 2835 54185
rect 2777 54145 2789 54179
rect 2823 54176 2835 54179
rect 2866 54176 2872 54188
rect 2823 54148 2872 54176
rect 2823 54145 2835 54148
rect 2777 54139 2835 54145
rect 1688 54108 1716 54139
rect 2866 54136 2872 54148
rect 2924 54136 2930 54188
rect 2961 54179 3019 54185
rect 2961 54145 2973 54179
rect 3007 54176 3019 54179
rect 3510 54176 3516 54188
rect 3007 54148 3516 54176
rect 3007 54145 3019 54148
rect 2961 54139 3019 54145
rect 3510 54136 3516 54148
rect 3568 54136 3574 54188
rect 9858 54176 9864 54188
rect 9819 54148 9864 54176
rect 9858 54136 9864 54148
rect 9916 54136 9922 54188
rect 7098 54108 7104 54120
rect 1688 54080 7104 54108
rect 7098 54068 7104 54080
rect 7156 54068 7162 54120
rect 10042 54040 10048 54052
rect 10003 54012 10048 54040
rect 10042 54000 10048 54012
rect 10100 54000 10106 54052
rect 1486 53972 1492 53984
rect 1447 53944 1492 53972
rect 1486 53932 1492 53944
rect 1544 53932 1550 53984
rect 2961 53975 3019 53981
rect 2961 53941 2973 53975
rect 3007 53972 3019 53975
rect 9858 53972 9864 53984
rect 3007 53944 9864 53972
rect 3007 53941 3019 53944
rect 2961 53935 3019 53941
rect 9858 53932 9864 53944
rect 9916 53932 9922 53984
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5845 53882
rect 5897 53830 5909 53882
rect 5961 53830 5973 53882
rect 6025 53830 6037 53882
rect 6089 53830 6101 53882
rect 6153 53830 9109 53882
rect 9161 53830 9173 53882
rect 9225 53830 9237 53882
rect 9289 53830 9301 53882
rect 9353 53830 9365 53882
rect 9417 53830 10856 53882
rect 1104 53808 10856 53830
rect 1578 53728 1584 53780
rect 1636 53768 1642 53780
rect 1636 53740 1900 53768
rect 1636 53728 1642 53740
rect 1762 53660 1768 53712
rect 1820 53660 1826 53712
rect 1780 53632 1808 53660
rect 1596 53604 1808 53632
rect 753 53567 811 53573
rect 753 53533 765 53567
rect 799 53564 811 53567
rect 1302 53564 1308 53576
rect 799 53536 1308 53564
rect 799 53533 811 53536
rect 753 53527 811 53533
rect 1302 53524 1308 53536
rect 1360 53564 1366 53576
rect 1596 53573 1624 53604
rect 1872 53573 1900 53740
rect 1946 53728 1952 53780
rect 2004 53768 2010 53780
rect 2685 53771 2743 53777
rect 2685 53768 2697 53771
rect 2004 53740 2697 53768
rect 2004 53728 2010 53740
rect 2685 53737 2697 53740
rect 2731 53737 2743 53771
rect 2685 53731 2743 53737
rect 8662 53700 8668 53712
rect 2240 53672 8668 53700
rect 1966 53635 2024 53641
rect 1966 53601 1978 53635
rect 2012 53632 2024 53635
rect 2240 53632 2268 53672
rect 8662 53660 8668 53672
rect 8720 53660 8726 53712
rect 2012 53604 2268 53632
rect 2012 53601 2024 53604
rect 1966 53595 2024 53601
rect 1397 53567 1455 53573
rect 1397 53564 1409 53567
rect 1360 53536 1409 53564
rect 1360 53524 1366 53536
rect 1397 53533 1409 53536
rect 1443 53533 1455 53567
rect 1397 53527 1455 53533
rect 1581 53567 1639 53573
rect 1581 53533 1593 53567
rect 1627 53533 1639 53567
rect 1581 53527 1639 53533
rect 1817 53567 1900 53573
rect 1817 53533 1829 53567
rect 1863 53536 1900 53567
rect 2501 53567 2559 53573
rect 1863 53533 1875 53536
rect 1817 53527 1875 53533
rect 2501 53533 2513 53567
rect 2547 53564 2559 53567
rect 2685 53567 2743 53573
rect 2547 53536 2636 53564
rect 2547 53533 2559 53536
rect 2501 53527 2559 53533
rect 2608 53508 2636 53536
rect 2685 53533 2697 53567
rect 2731 53564 2743 53567
rect 3326 53564 3332 53576
rect 2731 53536 3332 53564
rect 2731 53533 2743 53536
rect 2685 53527 2743 53533
rect 3326 53524 3332 53536
rect 3384 53524 3390 53576
rect 9861 53567 9919 53573
rect 9861 53533 9873 53567
rect 9907 53564 9919 53567
rect 11057 53567 11115 53573
rect 11057 53564 11069 53567
rect 9907 53536 11069 53564
rect 9907 53533 9919 53536
rect 9861 53527 9919 53533
rect 11057 53533 11069 53536
rect 11103 53533 11115 53567
rect 11057 53527 11115 53533
rect 1673 53499 1731 53505
rect 1673 53465 1685 53499
rect 1719 53496 1731 53499
rect 1719 53468 2452 53496
rect 1719 53465 1731 53468
rect 1673 53459 1731 53465
rect 845 53431 903 53437
rect 845 53397 857 53431
rect 891 53428 903 53431
rect 1854 53428 1860 53440
rect 891 53400 1860 53428
rect 891 53397 903 53400
rect 845 53391 903 53397
rect 1854 53388 1860 53400
rect 1912 53388 1918 53440
rect 2424 53428 2452 53468
rect 2590 53456 2596 53508
rect 2648 53496 2654 53508
rect 2958 53496 2964 53508
rect 2648 53468 2964 53496
rect 2648 53456 2654 53468
rect 2958 53456 2964 53468
rect 3016 53456 3022 53508
rect 9950 53496 9956 53508
rect 6288 53468 9956 53496
rect 6288 53428 6316 53468
rect 9950 53456 9956 53468
rect 10008 53456 10014 53508
rect 10042 53428 10048 53440
rect 2424 53400 6316 53428
rect 10003 53400 10048 53428
rect 10042 53388 10048 53400
rect 10100 53388 10106 53440
rect 11057 53431 11115 53437
rect 11057 53397 11069 53431
rect 11103 53428 11115 53431
rect 11333 53431 11391 53437
rect 11333 53428 11345 53431
rect 11103 53400 11345 53428
rect 11103 53397 11115 53400
rect 11057 53391 11115 53397
rect 11333 53397 11345 53400
rect 11379 53397 11391 53431
rect 11333 53391 11391 53397
rect 1104 53338 10856 53360
rect 1104 53286 4213 53338
rect 4265 53286 4277 53338
rect 4329 53286 4341 53338
rect 4393 53286 4405 53338
rect 4457 53286 4469 53338
rect 4521 53286 7477 53338
rect 7529 53286 7541 53338
rect 7593 53286 7605 53338
rect 7657 53286 7669 53338
rect 7721 53286 7733 53338
rect 7785 53286 10856 53338
rect 1104 53264 10856 53286
rect 2424 53196 2636 53224
rect 2424 53156 2452 53196
rect 1688 53128 2452 53156
rect 2608 53156 2636 53196
rect 7282 53156 7288 53168
rect 2608 53128 7288 53156
rect 1688 53097 1716 53128
rect 7282 53116 7288 53128
rect 7340 53116 7346 53168
rect 1673 53091 1731 53097
rect 1673 53057 1685 53091
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 1946 53048 1952 53100
rect 2004 53088 2010 53100
rect 2133 53091 2191 53097
rect 2133 53088 2145 53091
rect 2004 53060 2145 53088
rect 2004 53048 2010 53060
rect 2133 53057 2145 53060
rect 2179 53057 2191 53091
rect 2133 53051 2191 53057
rect 2869 53091 2927 53097
rect 2869 53057 2881 53091
rect 2915 53088 2927 53091
rect 7374 53088 7380 53100
rect 2915 53060 7380 53088
rect 2915 53057 2927 53060
rect 2869 53051 2927 53057
rect 7374 53048 7380 53060
rect 7432 53048 7438 53100
rect 9858 53088 9864 53100
rect 9819 53060 9864 53088
rect 9858 53048 9864 53060
rect 9916 53048 9922 53100
rect 290 52912 296 52964
rect 348 52952 354 52964
rect 2590 52952 2596 52964
rect 348 52924 2596 52952
rect 348 52912 354 52924
rect 2590 52912 2596 52924
rect 2648 52912 2654 52964
rect 3050 52952 3056 52964
rect 3011 52924 3056 52952
rect 3050 52912 3056 52924
rect 3108 52912 3114 52964
rect 1394 52844 1400 52896
rect 1452 52884 1458 52896
rect 1489 52887 1547 52893
rect 1489 52884 1501 52887
rect 1452 52856 1501 52884
rect 1452 52844 1458 52856
rect 1489 52853 1501 52856
rect 1535 52853 1547 52887
rect 2314 52884 2320 52896
rect 2275 52856 2320 52884
rect 1489 52847 1547 52853
rect 2314 52844 2320 52856
rect 2372 52844 2378 52896
rect 10042 52884 10048 52896
rect 10003 52856 10048 52884
rect 10042 52844 10048 52856
rect 10100 52844 10106 52896
rect 1104 52794 10856 52816
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5845 52794
rect 5897 52742 5909 52794
rect 5961 52742 5973 52794
rect 6025 52742 6037 52794
rect 6089 52742 6101 52794
rect 6153 52742 9109 52794
rect 9161 52742 9173 52794
rect 9225 52742 9237 52794
rect 9289 52742 9301 52794
rect 9353 52742 9365 52794
rect 9417 52742 10856 52794
rect 1104 52720 10856 52742
rect 1946 52640 1952 52692
rect 2004 52640 2010 52692
rect 2222 52680 2228 52692
rect 2183 52652 2228 52680
rect 2222 52640 2228 52652
rect 2280 52640 2286 52692
rect 1964 52612 1992 52640
rect 6270 52612 6276 52624
rect 1964 52584 6276 52612
rect 6270 52572 6276 52584
rect 6328 52572 6334 52624
rect 2590 52544 2596 52556
rect 2240 52516 2596 52544
rect 1673 52479 1731 52485
rect 1673 52445 1685 52479
rect 1719 52476 1731 52479
rect 1854 52476 1860 52488
rect 1719 52448 1860 52476
rect 1719 52445 1731 52448
rect 1673 52439 1731 52445
rect 1854 52436 1860 52448
rect 1912 52436 1918 52488
rect 2240 52485 2268 52516
rect 2590 52504 2596 52516
rect 2648 52544 2654 52556
rect 3326 52544 3332 52556
rect 2648 52516 3332 52544
rect 2648 52504 2654 52516
rect 3326 52504 3332 52516
rect 3384 52504 3390 52556
rect 2225 52479 2283 52485
rect 2225 52445 2237 52479
rect 2271 52445 2283 52479
rect 2225 52439 2283 52445
rect 2314 52436 2320 52488
rect 2372 52476 2378 52488
rect 2409 52479 2467 52485
rect 2409 52476 2421 52479
rect 2372 52448 2421 52476
rect 2372 52436 2378 52448
rect 2409 52445 2421 52448
rect 2455 52445 2467 52479
rect 2409 52439 2467 52445
rect 1486 52340 1492 52352
rect 1447 52312 1492 52340
rect 1486 52300 1492 52312
rect 1544 52300 1550 52352
rect 1104 52250 10856 52272
rect 1104 52198 4213 52250
rect 4265 52198 4277 52250
rect 4329 52198 4341 52250
rect 4393 52198 4405 52250
rect 4457 52198 4469 52250
rect 4521 52198 7477 52250
rect 7529 52198 7541 52250
rect 7593 52198 7605 52250
rect 7657 52198 7669 52250
rect 7721 52198 7733 52250
rect 7785 52198 10856 52250
rect 1104 52176 10856 52198
rect 1762 52136 1768 52148
rect 1596 52108 1768 52136
rect 1596 52077 1624 52108
rect 1762 52096 1768 52108
rect 1820 52096 1826 52148
rect 1946 52096 1952 52148
rect 2004 52136 2010 52148
rect 2501 52139 2559 52145
rect 2501 52136 2513 52139
rect 2004 52108 2513 52136
rect 2004 52096 2010 52108
rect 2501 52105 2513 52108
rect 2547 52105 2559 52139
rect 2501 52099 2559 52105
rect 1581 52071 1639 52077
rect 1581 52037 1593 52071
rect 1627 52037 1639 52071
rect 1581 52031 1639 52037
rect 1673 52071 1731 52077
rect 1673 52037 1685 52071
rect 1719 52068 1731 52071
rect 11241 52071 11299 52077
rect 11241 52068 11253 52071
rect 1719 52040 11253 52068
rect 1719 52037 1731 52040
rect 1673 52031 1731 52037
rect 11241 52037 11253 52040
rect 11287 52037 11299 52071
rect 11241 52031 11299 52037
rect 1302 51960 1308 52012
rect 1360 52000 1366 52012
rect 1397 52003 1455 52009
rect 1397 52000 1409 52003
rect 1360 51972 1409 52000
rect 1360 51960 1366 51972
rect 1397 51969 1409 51972
rect 1443 51969 1455 52003
rect 1397 51963 1455 51969
rect 1765 52003 1823 52009
rect 1765 51969 1777 52003
rect 1811 51969 1823 52003
rect 1765 51963 1823 51969
rect 2409 52003 2467 52009
rect 2409 51969 2421 52003
rect 2455 52000 2467 52003
rect 2590 52000 2596 52012
rect 2455 51972 2489 52000
rect 2551 51972 2596 52000
rect 2455 51969 2467 51972
rect 2409 51963 2467 51969
rect 1578 51824 1584 51876
rect 1636 51864 1642 51876
rect 1780 51864 1808 51963
rect 2424 51932 2452 51963
rect 2590 51960 2596 51972
rect 2648 52000 2654 52012
rect 2958 52000 2964 52012
rect 2648 51972 2964 52000
rect 2648 51960 2654 51972
rect 2958 51960 2964 51972
rect 3016 51960 3022 52012
rect 3053 52003 3111 52009
rect 3053 51969 3065 52003
rect 3099 51969 3111 52003
rect 3053 51963 3111 51969
rect 3237 52003 3295 52009
rect 3237 51969 3249 52003
rect 3283 52000 3295 52003
rect 3510 52000 3516 52012
rect 3283 51972 3516 52000
rect 3283 51969 3295 51972
rect 3237 51963 3295 51969
rect 3068 51932 3096 51963
rect 3510 51960 3516 51972
rect 3568 51960 3574 52012
rect 9861 52003 9919 52009
rect 9861 51969 9873 52003
rect 9907 51969 9919 52003
rect 9861 51963 9919 51969
rect 1636 51836 1808 51864
rect 1872 51904 3096 51932
rect 3145 51935 3203 51941
rect 1636 51824 1642 51836
rect 474 51756 480 51808
rect 532 51796 538 51808
rect 1872 51796 1900 51904
rect 3145 51901 3157 51935
rect 3191 51932 3203 51935
rect 9876 51932 9904 51963
rect 3191 51904 9904 51932
rect 11241 51935 11299 51941
rect 3191 51901 3203 51904
rect 3145 51895 3203 51901
rect 11241 51901 11253 51935
rect 11287 51932 11299 51935
rect 11885 51935 11943 51941
rect 11885 51932 11897 51935
rect 11287 51904 11897 51932
rect 11287 51901 11299 51904
rect 11241 51895 11299 51901
rect 11885 51901 11897 51904
rect 11931 51901 11943 51935
rect 11885 51895 11943 51901
rect 1949 51867 2007 51873
rect 1949 51833 1961 51867
rect 1995 51864 2007 51867
rect 3326 51864 3332 51876
rect 1995 51836 3332 51864
rect 1995 51833 2007 51836
rect 1949 51827 2007 51833
rect 3326 51824 3332 51836
rect 3384 51824 3390 51876
rect 10042 51796 10048 51808
rect 532 51768 1900 51796
rect 10003 51768 10048 51796
rect 532 51756 538 51768
rect 10042 51756 10048 51768
rect 10100 51756 10106 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5845 51706
rect 5897 51654 5909 51706
rect 5961 51654 5973 51706
rect 6025 51654 6037 51706
rect 6089 51654 6101 51706
rect 6153 51654 9109 51706
rect 9161 51654 9173 51706
rect 9225 51654 9237 51706
rect 9289 51654 9301 51706
rect 9353 51654 9365 51706
rect 9417 51654 10856 51706
rect 1104 51632 10856 51654
rect 7926 51456 7932 51468
rect 1688 51428 7932 51456
rect 1688 51397 1716 51428
rect 7926 51416 7932 51428
rect 7984 51416 7990 51468
rect 1673 51391 1731 51397
rect 1673 51357 1685 51391
rect 1719 51357 1731 51391
rect 1673 51351 1731 51357
rect 2409 51391 2467 51397
rect 2409 51357 2421 51391
rect 2455 51357 2467 51391
rect 2409 51351 2467 51357
rect 2424 51320 2452 51351
rect 2774 51348 2780 51400
rect 2832 51388 2838 51400
rect 2869 51391 2927 51397
rect 2869 51388 2881 51391
rect 2832 51360 2881 51388
rect 2832 51348 2838 51360
rect 2869 51357 2881 51360
rect 2915 51357 2927 51391
rect 9858 51388 9864 51400
rect 9819 51360 9864 51388
rect 2869 51351 2927 51357
rect 9858 51348 9864 51360
rect 9916 51348 9922 51400
rect 7834 51320 7840 51332
rect 2424 51292 7840 51320
rect 7834 51280 7840 51292
rect 7892 51280 7898 51332
rect 1394 51212 1400 51264
rect 1452 51252 1458 51264
rect 1489 51255 1547 51261
rect 1489 51252 1501 51255
rect 1452 51224 1501 51252
rect 1452 51212 1458 51224
rect 1489 51221 1501 51224
rect 1535 51221 1547 51255
rect 2222 51252 2228 51264
rect 2183 51224 2228 51252
rect 1489 51215 1547 51221
rect 2222 51212 2228 51224
rect 2280 51212 2286 51264
rect 3050 51252 3056 51264
rect 3011 51224 3056 51252
rect 3050 51212 3056 51224
rect 3108 51212 3114 51264
rect 10042 51252 10048 51264
rect 10003 51224 10048 51252
rect 10042 51212 10048 51224
rect 10100 51212 10106 51264
rect 1104 51162 10856 51184
rect 1104 51110 4213 51162
rect 4265 51110 4277 51162
rect 4329 51110 4341 51162
rect 4393 51110 4405 51162
rect 4457 51110 4469 51162
rect 4521 51110 7477 51162
rect 7529 51110 7541 51162
rect 7593 51110 7605 51162
rect 7657 51110 7669 51162
rect 7721 51110 7733 51162
rect 7785 51110 10856 51162
rect 1104 51088 10856 51110
rect 3145 51051 3203 51057
rect 3145 51017 3157 51051
rect 3191 51048 3203 51051
rect 9858 51048 9864 51060
rect 3191 51020 9864 51048
rect 3191 51017 3203 51020
rect 3145 51011 3203 51017
rect 9858 51008 9864 51020
rect 9916 51008 9922 51060
rect 3510 50980 3516 50992
rect 3068 50952 3516 50980
rect 3068 50921 3096 50952
rect 3510 50940 3516 50952
rect 3568 50940 3574 50992
rect 1673 50915 1731 50921
rect 1673 50881 1685 50915
rect 1719 50912 1731 50915
rect 3053 50915 3111 50921
rect 1719 50884 2774 50912
rect 1719 50881 1731 50884
rect 1673 50875 1731 50881
rect 2746 50844 2774 50884
rect 3053 50881 3065 50915
rect 3099 50881 3111 50915
rect 3053 50875 3111 50881
rect 3237 50915 3295 50921
rect 3237 50881 3249 50915
rect 3283 50912 3295 50915
rect 4154 50912 4160 50924
rect 3283 50884 4160 50912
rect 3283 50881 3295 50884
rect 3237 50875 3295 50881
rect 4154 50872 4160 50884
rect 4212 50872 4218 50924
rect 7190 50844 7196 50856
rect 2746 50816 7196 50844
rect 7190 50804 7196 50816
rect 7248 50804 7254 50856
rect 2774 50736 2780 50788
rect 2832 50776 2838 50788
rect 3786 50776 3792 50788
rect 2832 50748 3792 50776
rect 2832 50736 2838 50748
rect 3786 50736 3792 50748
rect 3844 50736 3850 50788
rect 1486 50708 1492 50720
rect 1447 50680 1492 50708
rect 1486 50668 1492 50680
rect 1544 50668 1550 50720
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5845 50618
rect 5897 50566 5909 50618
rect 5961 50566 5973 50618
rect 6025 50566 6037 50618
rect 6089 50566 6101 50618
rect 6153 50566 9109 50618
rect 9161 50566 9173 50618
rect 9225 50566 9237 50618
rect 9289 50566 9301 50618
rect 9353 50566 9365 50618
rect 9417 50566 10856 50618
rect 1104 50544 10856 50566
rect 1302 50464 1308 50516
rect 1360 50504 1366 50516
rect 1946 50504 1952 50516
rect 1360 50476 1952 50504
rect 1360 50464 1366 50476
rect 1946 50464 1952 50476
rect 2004 50464 2010 50516
rect 2498 50464 2504 50516
rect 2556 50504 2562 50516
rect 2593 50507 2651 50513
rect 2593 50504 2605 50507
rect 2556 50476 2605 50504
rect 2556 50464 2562 50476
rect 2593 50473 2605 50476
rect 2639 50473 2651 50507
rect 2593 50467 2651 50473
rect 3053 50507 3111 50513
rect 3053 50473 3065 50507
rect 3099 50504 3111 50507
rect 3694 50504 3700 50516
rect 3099 50476 3700 50504
rect 3099 50473 3111 50476
rect 3053 50467 3111 50473
rect 3694 50464 3700 50476
rect 3752 50464 3758 50516
rect 3973 50507 4031 50513
rect 3973 50473 3985 50507
rect 4019 50504 4031 50507
rect 4019 50476 9904 50504
rect 4019 50473 4031 50476
rect 3973 50467 4031 50473
rect 1670 50396 1676 50448
rect 1728 50436 1734 50448
rect 2406 50436 2412 50448
rect 1728 50408 2412 50436
rect 1728 50396 1734 50408
rect 2406 50396 2412 50408
rect 2464 50396 2470 50448
rect 3510 50396 3516 50448
rect 3568 50436 3574 50448
rect 3568 50408 3924 50436
rect 3568 50396 3574 50408
rect 1302 50328 1308 50380
rect 1360 50368 1366 50380
rect 1360 50340 3832 50368
rect 1360 50328 1366 50340
rect 1578 50300 1584 50312
rect 1539 50272 1584 50300
rect 1578 50260 1584 50272
rect 1636 50260 1642 50312
rect 1673 50303 1731 50309
rect 1673 50269 1685 50303
rect 1719 50300 1731 50303
rect 1719 50272 1900 50300
rect 1719 50269 1731 50272
rect 1673 50263 1731 50269
rect 1026 50192 1032 50244
rect 1084 50232 1090 50244
rect 1765 50235 1823 50241
rect 1765 50232 1777 50235
rect 1084 50204 1777 50232
rect 1084 50192 1090 50204
rect 1765 50201 1777 50204
rect 1811 50201 1823 50235
rect 1872 50232 1900 50272
rect 1946 50260 1952 50312
rect 2004 50300 2010 50312
rect 2424 50309 2452 50340
rect 2409 50303 2467 50309
rect 2004 50272 2049 50300
rect 2004 50260 2010 50272
rect 2409 50269 2421 50303
rect 2455 50269 2467 50303
rect 2409 50263 2467 50269
rect 2593 50303 2651 50309
rect 2593 50269 2605 50303
rect 2639 50300 2651 50303
rect 2958 50300 2964 50312
rect 2639 50272 2964 50300
rect 2639 50269 2651 50272
rect 2593 50263 2651 50269
rect 2958 50260 2964 50272
rect 3016 50300 3022 50312
rect 3804 50309 3832 50340
rect 3053 50303 3111 50309
rect 3053 50300 3065 50303
rect 3016 50272 3065 50300
rect 3016 50260 3022 50272
rect 3053 50269 3065 50272
rect 3099 50269 3111 50303
rect 3053 50263 3111 50269
rect 3237 50303 3295 50309
rect 3237 50269 3249 50303
rect 3283 50269 3295 50303
rect 3237 50263 3295 50269
rect 3789 50303 3847 50309
rect 3789 50269 3801 50303
rect 3835 50269 3847 50303
rect 3896 50300 3924 50408
rect 9876 50309 9904 50476
rect 3973 50303 4031 50309
rect 3973 50300 3985 50303
rect 3896 50272 3985 50300
rect 3789 50263 3847 50269
rect 3973 50269 3985 50272
rect 4019 50269 4031 50303
rect 3973 50263 4031 50269
rect 9861 50303 9919 50309
rect 9861 50269 9873 50303
rect 9907 50269 9919 50303
rect 9861 50263 9919 50269
rect 3252 50232 3280 50263
rect 4154 50232 4160 50244
rect 1872 50204 2774 50232
rect 3252 50204 4160 50232
rect 1765 50195 1823 50201
rect 1397 50167 1455 50173
rect 1397 50133 1409 50167
rect 1443 50164 1455 50167
rect 1670 50164 1676 50176
rect 1443 50136 1676 50164
rect 1443 50133 1455 50136
rect 1397 50127 1455 50133
rect 1670 50124 1676 50136
rect 1728 50124 1734 50176
rect 2746 50164 2774 50204
rect 4154 50192 4160 50204
rect 4212 50232 4218 50244
rect 4614 50232 4620 50244
rect 4212 50204 4620 50232
rect 4212 50192 4218 50204
rect 4614 50192 4620 50204
rect 4672 50192 4678 50244
rect 11793 50235 11851 50241
rect 11793 50232 11805 50235
rect 4724 50204 11805 50232
rect 4724 50164 4752 50204
rect 11793 50201 11805 50204
rect 11839 50201 11851 50235
rect 11793 50195 11851 50201
rect 10042 50164 10048 50176
rect 2746 50136 4752 50164
rect 10003 50136 10048 50164
rect 10042 50124 10048 50136
rect 10100 50124 10106 50176
rect 1104 50074 10856 50096
rect 1104 50022 4213 50074
rect 4265 50022 4277 50074
rect 4329 50022 4341 50074
rect 4393 50022 4405 50074
rect 4457 50022 4469 50074
rect 4521 50022 7477 50074
rect 7529 50022 7541 50074
rect 7593 50022 7605 50074
rect 7657 50022 7669 50074
rect 7721 50022 7733 50074
rect 7785 50022 10856 50074
rect 1104 50000 10856 50022
rect 1673 49895 1731 49901
rect 1673 49861 1685 49895
rect 1719 49892 1731 49895
rect 11609 49895 11667 49901
rect 11609 49892 11621 49895
rect 1719 49864 11621 49892
rect 1719 49861 1731 49864
rect 1673 49855 1731 49861
rect 11609 49861 11621 49864
rect 11655 49861 11667 49895
rect 11609 49855 11667 49861
rect 1578 49824 1584 49836
rect 1539 49796 1584 49824
rect 1578 49784 1584 49796
rect 1636 49784 1642 49836
rect 1765 49827 1823 49833
rect 1765 49793 1777 49827
rect 1811 49793 1823 49827
rect 1946 49824 1952 49836
rect 1907 49796 1952 49824
rect 1765 49787 1823 49793
rect 1118 49716 1124 49768
rect 1176 49756 1182 49768
rect 1780 49756 1808 49787
rect 1946 49784 1952 49796
rect 2004 49784 2010 49836
rect 2409 49827 2467 49833
rect 2409 49793 2421 49827
rect 2455 49824 2467 49827
rect 6178 49824 6184 49836
rect 2455 49796 6184 49824
rect 2455 49793 2467 49796
rect 2409 49787 2467 49793
rect 6178 49784 6184 49796
rect 6236 49784 6242 49836
rect 9858 49824 9864 49836
rect 9819 49796 9864 49824
rect 9858 49784 9864 49796
rect 9916 49784 9922 49836
rect 1176 49728 1808 49756
rect 1176 49716 1182 49728
rect 1486 49648 1492 49700
rect 1544 49688 1550 49700
rect 1964 49688 1992 49784
rect 3970 49716 3976 49768
rect 4028 49756 4034 49768
rect 5166 49756 5172 49768
rect 4028 49728 5172 49756
rect 4028 49716 4034 49728
rect 5166 49716 5172 49728
rect 5224 49716 5230 49768
rect 1544 49660 1992 49688
rect 1544 49648 1550 49660
rect 1394 49620 1400 49632
rect 1355 49592 1400 49620
rect 1394 49580 1400 49592
rect 1452 49580 1458 49632
rect 1946 49580 1952 49632
rect 2004 49620 2010 49632
rect 2314 49620 2320 49632
rect 2004 49592 2320 49620
rect 2004 49580 2010 49592
rect 2314 49580 2320 49592
rect 2372 49580 2378 49632
rect 2406 49580 2412 49632
rect 2464 49620 2470 49632
rect 2593 49623 2651 49629
rect 2593 49620 2605 49623
rect 2464 49592 2605 49620
rect 2464 49580 2470 49592
rect 2593 49589 2605 49592
rect 2639 49589 2651 49623
rect 2593 49583 2651 49589
rect 4614 49580 4620 49632
rect 4672 49620 4678 49632
rect 5166 49620 5172 49632
rect 4672 49592 5172 49620
rect 4672 49580 4678 49592
rect 5166 49580 5172 49592
rect 5224 49580 5230 49632
rect 10042 49620 10048 49632
rect 10003 49592 10048 49620
rect 10042 49580 10048 49592
rect 10100 49580 10106 49632
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5845 49530
rect 5897 49478 5909 49530
rect 5961 49478 5973 49530
rect 6025 49478 6037 49530
rect 6089 49478 6101 49530
rect 6153 49478 9109 49530
rect 9161 49478 9173 49530
rect 9225 49478 9237 49530
rect 9289 49478 9301 49530
rect 9353 49478 9365 49530
rect 9417 49478 10856 49530
rect 1104 49456 10856 49478
rect 11701 49419 11759 49425
rect 11701 49416 11713 49419
rect 1688 49388 11713 49416
rect 1397 49215 1455 49221
rect 1397 49181 1409 49215
rect 1443 49212 1455 49215
rect 1486 49212 1492 49224
rect 1443 49184 1492 49212
rect 1443 49181 1455 49184
rect 1397 49175 1455 49181
rect 1486 49172 1492 49184
rect 1544 49172 1550 49224
rect 1688 49221 1716 49388
rect 11701 49385 11713 49388
rect 11747 49385 11759 49419
rect 11701 49379 11759 49385
rect 6730 49280 6736 49292
rect 2746 49252 6736 49280
rect 1673 49215 1731 49221
rect 1673 49181 1685 49215
rect 1719 49181 1731 49215
rect 1673 49175 1731 49181
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49181 1823 49215
rect 1765 49175 1823 49181
rect 2409 49215 2467 49221
rect 2409 49181 2421 49215
rect 2455 49212 2467 49215
rect 2746 49212 2774 49252
rect 6730 49240 6736 49252
rect 6788 49240 6794 49292
rect 2455 49184 2774 49212
rect 2455 49181 2467 49184
rect 2409 49175 2467 49181
rect 382 49104 388 49156
rect 440 49144 446 49156
rect 1581 49147 1639 49153
rect 1581 49144 1593 49147
rect 440 49116 1593 49144
rect 440 49104 446 49116
rect 1581 49113 1593 49116
rect 1627 49113 1639 49147
rect 1780 49144 1808 49175
rect 3510 49172 3516 49224
rect 3568 49212 3574 49224
rect 3789 49215 3847 49221
rect 3789 49212 3801 49215
rect 3568 49184 3801 49212
rect 3568 49172 3574 49184
rect 3789 49181 3801 49184
rect 3835 49212 3847 49215
rect 4614 49212 4620 49224
rect 3835 49184 4620 49212
rect 3835 49181 3847 49184
rect 3789 49175 3847 49181
rect 4614 49172 4620 49184
rect 4672 49172 4678 49224
rect 9766 49172 9772 49224
rect 9824 49212 9830 49224
rect 9861 49215 9919 49221
rect 9861 49212 9873 49215
rect 9824 49184 9873 49212
rect 9824 49172 9830 49184
rect 9861 49181 9873 49184
rect 9907 49181 9919 49215
rect 9861 49175 9919 49181
rect 4065 49147 4123 49153
rect 4065 49144 4077 49147
rect 1581 49107 1639 49113
rect 1688 49116 1808 49144
rect 3528 49116 4077 49144
rect 1486 49036 1492 49088
rect 1544 49076 1550 49088
rect 1688 49076 1716 49116
rect 3528 49088 3556 49116
rect 4065 49113 4077 49116
rect 4111 49113 4123 49147
rect 4065 49107 4123 49113
rect 1544 49048 1716 49076
rect 1949 49079 2007 49085
rect 1544 49036 1550 49048
rect 1949 49045 1961 49079
rect 1995 49076 2007 49079
rect 2314 49076 2320 49088
rect 1995 49048 2320 49076
rect 1995 49045 2007 49048
rect 1949 49039 2007 49045
rect 2314 49036 2320 49048
rect 2372 49036 2378 49088
rect 2593 49079 2651 49085
rect 2593 49045 2605 49079
rect 2639 49076 2651 49079
rect 2774 49076 2780 49088
rect 2639 49048 2780 49076
rect 2639 49045 2651 49048
rect 2593 49039 2651 49045
rect 2774 49036 2780 49048
rect 2832 49036 2838 49088
rect 3510 49036 3516 49088
rect 3568 49036 3574 49088
rect 10042 49076 10048 49088
rect 10003 49048 10048 49076
rect 10042 49036 10048 49048
rect 10100 49036 10106 49088
rect 1104 48986 10856 49008
rect 1104 48934 4213 48986
rect 4265 48934 4277 48986
rect 4329 48934 4341 48986
rect 4393 48934 4405 48986
rect 4457 48934 4469 48986
rect 4521 48934 7477 48986
rect 7529 48934 7541 48986
rect 7593 48934 7605 48986
rect 7657 48934 7669 48986
rect 7721 48934 7733 48986
rect 7785 48934 10856 48986
rect 1104 48912 10856 48934
rect 382 48832 388 48884
rect 440 48872 446 48884
rect 1302 48872 1308 48884
rect 440 48844 1308 48872
rect 440 48832 446 48844
rect 1302 48832 1308 48844
rect 1360 48832 1366 48884
rect 2222 48872 2228 48884
rect 2183 48844 2228 48872
rect 2222 48832 2228 48844
rect 2280 48832 2286 48884
rect 1673 48739 1731 48745
rect 1673 48705 1685 48739
rect 1719 48705 1731 48739
rect 1673 48699 1731 48705
rect 2409 48739 2467 48745
rect 2409 48705 2421 48739
rect 2455 48736 2467 48739
rect 6546 48736 6552 48748
rect 2455 48708 6552 48736
rect 2455 48705 2467 48708
rect 2409 48699 2467 48705
rect 1688 48668 1716 48699
rect 6546 48696 6552 48708
rect 6604 48696 6610 48748
rect 6454 48668 6460 48680
rect 1688 48640 6460 48668
rect 6454 48628 6460 48640
rect 6512 48628 6518 48680
rect 2222 48560 2228 48612
rect 2280 48600 2286 48612
rect 2406 48600 2412 48612
rect 2280 48572 2412 48600
rect 2280 48560 2286 48572
rect 2406 48560 2412 48572
rect 2464 48560 2470 48612
rect 1486 48532 1492 48544
rect 1447 48504 1492 48532
rect 1486 48492 1492 48504
rect 1544 48492 1550 48544
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5845 48442
rect 5897 48390 5909 48442
rect 5961 48390 5973 48442
rect 6025 48390 6037 48442
rect 6089 48390 6101 48442
rect 6153 48390 9109 48442
rect 9161 48390 9173 48442
rect 9225 48390 9237 48442
rect 9289 48390 9301 48442
rect 9353 48390 9365 48442
rect 9417 48390 10856 48442
rect 1104 48368 10856 48390
rect 14 48288 20 48340
rect 72 48328 78 48340
rect 1578 48328 1584 48340
rect 72 48300 1584 48328
rect 72 48288 78 48300
rect 1578 48288 1584 48300
rect 1636 48288 1642 48340
rect 2406 48288 2412 48340
rect 2464 48328 2470 48340
rect 5534 48328 5540 48340
rect 2464 48300 5540 48328
rect 2464 48288 2470 48300
rect 5534 48288 5540 48300
rect 5592 48288 5598 48340
rect 2866 48220 2872 48272
rect 2924 48260 2930 48272
rect 3050 48260 3056 48272
rect 2924 48232 3056 48260
rect 2924 48220 2930 48232
rect 3050 48220 3056 48232
rect 3108 48220 3114 48272
rect 753 48195 811 48201
rect 753 48161 765 48195
rect 799 48192 811 48195
rect 4522 48192 4528 48204
rect 799 48164 4528 48192
rect 799 48161 811 48164
rect 753 48155 811 48161
rect 4522 48152 4528 48164
rect 4580 48152 4586 48204
rect 1673 48127 1731 48133
rect 1673 48093 1685 48127
rect 1719 48093 1731 48127
rect 1673 48087 1731 48093
rect 1688 48056 1716 48087
rect 1946 48084 1952 48136
rect 2004 48124 2010 48136
rect 2593 48127 2651 48133
rect 2593 48124 2605 48127
rect 2004 48096 2605 48124
rect 2004 48084 2010 48096
rect 2593 48093 2605 48096
rect 2639 48093 2651 48127
rect 2774 48124 2780 48136
rect 2735 48096 2780 48124
rect 2593 48087 2651 48093
rect 2774 48084 2780 48096
rect 2832 48084 2838 48136
rect 3050 48084 3056 48136
rect 3108 48124 3114 48136
rect 9861 48127 9919 48133
rect 9861 48124 9873 48127
rect 3108 48096 9873 48124
rect 3108 48084 3114 48096
rect 9861 48093 9873 48096
rect 9907 48093 9919 48127
rect 9861 48087 9919 48093
rect 6178 48056 6184 48068
rect 1688 48028 6184 48056
rect 6178 48016 6184 48028
rect 6236 48016 6242 48068
rect 1486 47988 1492 48000
rect 1447 47960 1492 47988
rect 1486 47948 1492 47960
rect 1544 47948 1550 48000
rect 2685 47991 2743 47997
rect 2685 47957 2697 47991
rect 2731 47988 2743 47991
rect 9858 47988 9864 48000
rect 2731 47960 9864 47988
rect 2731 47957 2743 47960
rect 2685 47951 2743 47957
rect 9858 47948 9864 47960
rect 9916 47948 9922 48000
rect 10042 47988 10048 48000
rect 10003 47960 10048 47988
rect 10042 47948 10048 47960
rect 10100 47948 10106 48000
rect 1104 47898 10856 47920
rect 1104 47846 4213 47898
rect 4265 47846 4277 47898
rect 4329 47846 4341 47898
rect 4393 47846 4405 47898
rect 4457 47846 4469 47898
rect 4521 47846 7477 47898
rect 7529 47846 7541 47898
rect 7593 47846 7605 47898
rect 7657 47846 7669 47898
rect 7721 47846 7733 47898
rect 7785 47846 10856 47898
rect 1104 47824 10856 47846
rect 2958 47784 2964 47796
rect 2919 47756 2964 47784
rect 2958 47744 2964 47756
rect 3016 47744 3022 47796
rect 3510 47744 3516 47796
rect 3568 47744 3574 47796
rect 661 47719 719 47725
rect 661 47685 673 47719
rect 707 47716 719 47719
rect 2498 47716 2504 47728
rect 707 47688 2504 47716
rect 707 47685 719 47688
rect 661 47679 719 47685
rect 2498 47676 2504 47688
rect 2556 47676 2562 47728
rect 3528 47716 3556 47744
rect 3528 47688 3740 47716
rect 1302 47608 1308 47660
rect 1360 47648 1366 47660
rect 1673 47651 1731 47657
rect 1673 47648 1685 47651
rect 1360 47620 1685 47648
rect 1360 47608 1366 47620
rect 1673 47617 1685 47620
rect 1719 47617 1731 47651
rect 1673 47611 1731 47617
rect 2409 47651 2467 47657
rect 2409 47617 2421 47651
rect 2455 47648 2467 47651
rect 2682 47648 2688 47660
rect 2455 47620 2688 47648
rect 2455 47617 2467 47620
rect 2409 47611 2467 47617
rect 2682 47608 2688 47620
rect 2740 47608 2746 47660
rect 2866 47648 2872 47660
rect 2827 47620 2872 47648
rect 2866 47608 2872 47620
rect 2924 47608 2930 47660
rect 2958 47608 2964 47660
rect 3016 47648 3022 47660
rect 3053 47651 3111 47657
rect 3053 47648 3065 47651
rect 3016 47620 3065 47648
rect 3016 47608 3022 47620
rect 3053 47617 3065 47620
rect 3099 47617 3111 47651
rect 3510 47648 3516 47660
rect 3471 47620 3516 47648
rect 3053 47611 3111 47617
rect 3510 47608 3516 47620
rect 3568 47608 3574 47660
rect 3712 47657 3740 47688
rect 3697 47651 3755 47657
rect 3697 47617 3709 47651
rect 3743 47617 3755 47651
rect 3697 47611 3755 47617
rect 9861 47651 9919 47657
rect 9861 47617 9873 47651
rect 9907 47617 9919 47651
rect 9861 47611 9919 47617
rect 1486 47540 1492 47592
rect 1544 47580 1550 47592
rect 1544 47552 2268 47580
rect 1544 47540 1550 47552
rect 2130 47512 2136 47524
rect 1044 47484 2136 47512
rect 1044 47240 1072 47484
rect 2130 47472 2136 47484
rect 2188 47472 2194 47524
rect 2240 47521 2268 47552
rect 2498 47540 2504 47592
rect 2556 47580 2562 47592
rect 2884 47580 2912 47608
rect 2556 47552 2912 47580
rect 3605 47583 3663 47589
rect 2556 47540 2562 47552
rect 3605 47549 3617 47583
rect 3651 47580 3663 47583
rect 9876 47580 9904 47611
rect 3651 47552 9904 47580
rect 3651 47549 3663 47552
rect 3605 47543 3663 47549
rect 2225 47515 2283 47521
rect 2225 47481 2237 47515
rect 2271 47481 2283 47515
rect 2225 47475 2283 47481
rect 1486 47444 1492 47456
rect 1447 47416 1492 47444
rect 1486 47404 1492 47416
rect 1544 47404 1550 47456
rect 10042 47444 10048 47456
rect 10003 47416 10048 47444
rect 10042 47404 10048 47416
rect 10100 47404 10106 47456
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5845 47354
rect 5897 47302 5909 47354
rect 5961 47302 5973 47354
rect 6025 47302 6037 47354
rect 6089 47302 6101 47354
rect 6153 47302 9109 47354
rect 9161 47302 9173 47354
rect 9225 47302 9237 47354
rect 9289 47302 9301 47354
rect 9353 47302 9365 47354
rect 9417 47302 10856 47354
rect 1104 47280 10856 47302
rect 2409 47243 2467 47249
rect 2409 47240 2421 47243
rect 1044 47212 2421 47240
rect 2409 47209 2421 47212
rect 2455 47209 2467 47243
rect 3050 47240 3056 47252
rect 3011 47212 3056 47240
rect 2409 47203 2467 47209
rect 3050 47200 3056 47212
rect 3108 47200 3114 47252
rect 1946 47132 1952 47184
rect 2004 47172 2010 47184
rect 2222 47172 2228 47184
rect 2004 47144 2228 47172
rect 2004 47132 2010 47144
rect 2222 47132 2228 47144
rect 2280 47132 2286 47184
rect 3510 47172 3516 47184
rect 2332 47144 3516 47172
rect 1026 47064 1032 47116
rect 1084 47104 1090 47116
rect 2332 47104 2360 47144
rect 3510 47132 3516 47144
rect 3568 47132 3574 47184
rect 1084 47076 1808 47104
rect 1084 47064 1090 47076
rect 1673 47039 1731 47045
rect 1673 47036 1685 47039
rect 1596 47008 1685 47036
rect 1486 46900 1492 46912
rect 1447 46872 1492 46900
rect 1486 46860 1492 46872
rect 1544 46860 1550 46912
rect 1596 46900 1624 47008
rect 1673 47005 1685 47008
rect 1719 47005 1731 47039
rect 1780 47036 1808 47076
rect 2240 47076 2360 47104
rect 2240 47045 2268 47076
rect 2225 47039 2283 47045
rect 2225 47036 2237 47039
rect 1780 47008 2237 47036
rect 1673 46999 1731 47005
rect 2225 47005 2237 47008
rect 2271 47005 2283 47039
rect 2225 46999 2283 47005
rect 2409 47039 2467 47045
rect 2409 47005 2421 47039
rect 2455 47036 2467 47039
rect 2498 47036 2504 47048
rect 2455 47008 2504 47036
rect 2455 47005 2467 47008
rect 2409 46999 2467 47005
rect 2498 46996 2504 47008
rect 2556 46996 2562 47048
rect 2866 47036 2872 47048
rect 2827 47008 2872 47036
rect 2866 46996 2872 47008
rect 2924 46996 2930 47048
rect 3053 47039 3111 47045
rect 3053 47036 3065 47039
rect 2976 47008 3065 47036
rect 2590 46900 2596 46912
rect 1596 46872 2596 46900
rect 2590 46860 2596 46872
rect 2648 46860 2654 46912
rect 2774 46860 2780 46912
rect 2832 46900 2838 46912
rect 2976 46900 3004 47008
rect 3053 47005 3065 47008
rect 3099 47005 3111 47039
rect 3053 46999 3111 47005
rect 2832 46872 3004 46900
rect 2832 46860 2838 46872
rect 1104 46810 10856 46832
rect 1104 46758 4213 46810
rect 4265 46758 4277 46810
rect 4329 46758 4341 46810
rect 4393 46758 4405 46810
rect 4457 46758 4469 46810
rect 4521 46758 7477 46810
rect 7529 46758 7541 46810
rect 7593 46758 7605 46810
rect 7657 46758 7669 46810
rect 7721 46758 7733 46810
rect 7785 46758 10856 46810
rect 1104 46736 10856 46758
rect 1118 46656 1124 46708
rect 1176 46696 1182 46708
rect 2866 46696 2872 46708
rect 1176 46668 2872 46696
rect 1176 46656 1182 46668
rect 2866 46656 2872 46668
rect 2924 46656 2930 46708
rect 10965 46699 11023 46705
rect 10965 46665 10977 46699
rect 11011 46696 11023 46699
rect 11333 46699 11391 46705
rect 11333 46696 11345 46699
rect 11011 46668 11345 46696
rect 11011 46665 11023 46668
rect 10965 46659 11023 46665
rect 11333 46665 11345 46668
rect 11379 46665 11391 46699
rect 11333 46659 11391 46665
rect 2590 46588 2596 46640
rect 2648 46628 2654 46640
rect 8938 46628 8944 46640
rect 2648 46600 8944 46628
rect 2648 46588 2654 46600
rect 8938 46588 8944 46600
rect 8996 46588 9002 46640
rect 1673 46563 1731 46569
rect 1673 46529 1685 46563
rect 1719 46529 1731 46563
rect 1673 46523 1731 46529
rect 1688 46492 1716 46523
rect 1946 46520 1952 46572
rect 2004 46560 2010 46572
rect 2501 46563 2559 46569
rect 2501 46560 2513 46563
rect 2004 46532 2513 46560
rect 2004 46520 2010 46532
rect 2501 46529 2513 46532
rect 2547 46529 2559 46563
rect 2501 46523 2559 46529
rect 2685 46563 2743 46569
rect 2685 46529 2697 46563
rect 2731 46560 2743 46563
rect 2774 46560 2780 46572
rect 2731 46532 2780 46560
rect 2731 46529 2743 46532
rect 2685 46523 2743 46529
rect 2774 46520 2780 46532
rect 2832 46520 2838 46572
rect 3510 46520 3516 46572
rect 3568 46560 3574 46572
rect 3786 46560 3792 46572
rect 3568 46532 3792 46560
rect 3568 46520 3574 46532
rect 3786 46520 3792 46532
rect 3844 46520 3850 46572
rect 9861 46563 9919 46569
rect 9861 46529 9873 46563
rect 9907 46560 9919 46563
rect 10965 46563 11023 46569
rect 10965 46560 10977 46563
rect 9907 46532 10977 46560
rect 9907 46529 9919 46532
rect 9861 46523 9919 46529
rect 10965 46529 10977 46532
rect 11011 46529 11023 46563
rect 10965 46523 11023 46529
rect 9030 46492 9036 46504
rect 1688 46464 9036 46492
rect 9030 46452 9036 46464
rect 9088 46452 9094 46504
rect 2685 46427 2743 46433
rect 2685 46393 2697 46427
rect 2731 46424 2743 46427
rect 9766 46424 9772 46436
rect 2731 46396 9772 46424
rect 2731 46393 2743 46396
rect 2685 46387 2743 46393
rect 9766 46384 9772 46396
rect 9824 46384 9830 46436
rect 10042 46424 10048 46436
rect 10003 46396 10048 46424
rect 10042 46384 10048 46396
rect 10100 46384 10106 46436
rect 1486 46356 1492 46368
rect 1447 46328 1492 46356
rect 1486 46316 1492 46328
rect 1544 46316 1550 46368
rect 4614 46316 4620 46368
rect 4672 46356 4678 46368
rect 5350 46356 5356 46368
rect 4672 46328 5356 46356
rect 4672 46316 4678 46328
rect 5350 46316 5356 46328
rect 5408 46316 5414 46368
rect 382 46288 388 46300
rect 124 46260 388 46288
rect 124 46096 152 46260
rect 382 46248 388 46260
rect 440 46248 446 46300
rect 1104 46266 10856 46288
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5845 46266
rect 5897 46214 5909 46266
rect 5961 46214 5973 46266
rect 6025 46214 6037 46266
rect 6089 46214 6101 46266
rect 6153 46214 9109 46266
rect 9161 46214 9173 46266
rect 9225 46214 9237 46266
rect 9289 46214 9301 46266
rect 9353 46214 9365 46266
rect 9417 46214 10856 46266
rect 1104 46192 10856 46214
rect 4798 46112 4804 46164
rect 4856 46152 4862 46164
rect 4982 46152 4988 46164
rect 4856 46124 4988 46152
rect 4856 46112 4862 46124
rect 4982 46112 4988 46124
rect 5040 46112 5046 46164
rect 106 46044 112 46096
rect 164 46044 170 46096
rect 474 46044 480 46096
rect 532 46084 538 46096
rect 1210 46084 1216 46096
rect 532 46056 1216 46084
rect 532 46044 538 46056
rect 1210 46044 1216 46056
rect 1268 46044 1274 46096
rect 3602 46044 3608 46096
rect 3660 46084 3666 46096
rect 4062 46084 4068 46096
rect 3660 46056 4068 46084
rect 3660 46044 3666 46056
rect 4062 46044 4068 46056
rect 4120 46044 4126 46096
rect 4522 46044 4528 46096
rect 4580 46084 4586 46096
rect 5350 46084 5356 46096
rect 4580 46056 5356 46084
rect 4580 46044 4586 46056
rect 5350 46044 5356 46056
rect 5408 46044 5414 46096
rect 4706 45976 4712 46028
rect 4764 46016 4770 46028
rect 4982 46016 4988 46028
rect 4764 45988 4988 46016
rect 4764 45976 4770 45988
rect 4982 45976 4988 45988
rect 5040 45976 5046 46028
rect 1673 45951 1731 45957
rect 1673 45917 1685 45951
rect 1719 45948 1731 45951
rect 8018 45948 8024 45960
rect 1719 45920 8024 45948
rect 1719 45917 1731 45920
rect 1673 45911 1731 45917
rect 8018 45908 8024 45920
rect 8076 45908 8082 45960
rect 9858 45948 9864 45960
rect 9819 45920 9864 45948
rect 9858 45908 9864 45920
rect 9916 45908 9922 45960
rect 4706 45840 4712 45892
rect 4764 45880 4770 45892
rect 5442 45880 5448 45892
rect 4764 45852 5448 45880
rect 4764 45840 4770 45852
rect 5442 45840 5448 45852
rect 5500 45840 5506 45892
rect 1486 45812 1492 45824
rect 1447 45784 1492 45812
rect 1486 45772 1492 45784
rect 1544 45772 1550 45824
rect 10042 45812 10048 45824
rect 10003 45784 10048 45812
rect 10042 45772 10048 45784
rect 10100 45772 10106 45824
rect 1104 45722 10856 45744
rect 1104 45670 4213 45722
rect 4265 45670 4277 45722
rect 4329 45670 4341 45722
rect 4393 45670 4405 45722
rect 4457 45670 4469 45722
rect 4521 45670 7477 45722
rect 7529 45670 7541 45722
rect 7593 45670 7605 45722
rect 7657 45670 7669 45722
rect 7721 45670 7733 45722
rect 7785 45670 10856 45722
rect 1104 45648 10856 45670
rect 1670 45568 1676 45620
rect 1728 45608 1734 45620
rect 1946 45608 1952 45620
rect 1728 45580 1952 45608
rect 1728 45568 1734 45580
rect 1946 45568 1952 45580
rect 2004 45568 2010 45620
rect 5166 45568 5172 45620
rect 5224 45608 5230 45620
rect 5350 45608 5356 45620
rect 5224 45580 5356 45608
rect 5224 45568 5230 45580
rect 5350 45568 5356 45580
rect 5408 45568 5414 45620
rect 845 45543 903 45549
rect 845 45509 857 45543
rect 891 45540 903 45543
rect 3418 45540 3424 45552
rect 891 45512 3424 45540
rect 891 45509 903 45512
rect 845 45503 903 45509
rect 3418 45500 3424 45512
rect 3476 45500 3482 45552
rect 1673 45475 1731 45481
rect 1673 45441 1685 45475
rect 1719 45441 1731 45475
rect 1673 45435 1731 45441
rect 1688 45336 1716 45435
rect 1946 45432 1952 45484
rect 2004 45472 2010 45484
rect 2317 45475 2375 45481
rect 2317 45472 2329 45475
rect 2004 45444 2329 45472
rect 2004 45432 2010 45444
rect 2317 45441 2329 45444
rect 2363 45441 2375 45475
rect 2317 45435 2375 45441
rect 1688 45308 2268 45336
rect 1486 45268 1492 45280
rect 1447 45240 1492 45268
rect 1486 45228 1492 45240
rect 1544 45228 1550 45280
rect 1854 45228 1860 45280
rect 1912 45268 1918 45280
rect 2133 45271 2191 45277
rect 2133 45268 2145 45271
rect 1912 45240 2145 45268
rect 1912 45228 1918 45240
rect 2133 45237 2145 45240
rect 2179 45237 2191 45271
rect 2240 45268 2268 45308
rect 5626 45268 5632 45280
rect 2240 45240 5632 45268
rect 2133 45231 2191 45237
rect 5626 45228 5632 45240
rect 5684 45228 5690 45280
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5845 45178
rect 5897 45126 5909 45178
rect 5961 45126 5973 45178
rect 6025 45126 6037 45178
rect 6089 45126 6101 45178
rect 6153 45126 9109 45178
rect 9161 45126 9173 45178
rect 9225 45126 9237 45178
rect 9289 45126 9301 45178
rect 9353 45126 9365 45178
rect 9417 45126 10856 45178
rect 1104 45104 10856 45126
rect 1486 45024 1492 45076
rect 1544 45064 1550 45076
rect 1544 45036 2774 45064
rect 1544 45024 1550 45036
rect 2746 45008 2774 45036
rect 4062 45024 4068 45076
rect 4120 45064 4126 45076
rect 5074 45064 5080 45076
rect 4120 45036 5080 45064
rect 4120 45024 4126 45036
rect 5074 45024 5080 45036
rect 5132 45024 5138 45076
rect 1762 44956 1768 45008
rect 1820 44996 1826 45008
rect 1949 44999 2007 45005
rect 1949 44996 1961 44999
rect 1820 44968 1961 44996
rect 1820 44956 1826 44968
rect 1949 44965 1961 44968
rect 1995 44965 2007 44999
rect 1949 44959 2007 44965
rect 2498 44956 2504 45008
rect 2556 44956 2562 45008
rect 2746 44968 2780 45008
rect 2774 44956 2780 44968
rect 2832 44956 2838 45008
rect 2222 44928 2228 44940
rect 1780 44900 2228 44928
rect 1780 44869 1808 44900
rect 2222 44888 2228 44900
rect 2280 44888 2286 44940
rect 2516 44928 2544 44956
rect 2332 44900 2544 44928
rect 1765 44863 1823 44869
rect 1765 44829 1777 44863
rect 1811 44829 1823 44863
rect 1765 44823 1823 44829
rect 1949 44863 2007 44869
rect 1949 44829 1961 44863
rect 1995 44860 2007 44863
rect 2332 44860 2360 44900
rect 1995 44832 2360 44860
rect 2501 44863 2559 44869
rect 1995 44829 2007 44832
rect 1949 44823 2007 44829
rect 2501 44829 2513 44863
rect 2547 44860 2559 44863
rect 6822 44860 6828 44872
rect 2547 44832 6828 44860
rect 2547 44829 2559 44832
rect 2501 44823 2559 44829
rect 6822 44820 6828 44832
rect 6880 44820 6886 44872
rect 9674 44820 9680 44872
rect 9732 44860 9738 44872
rect 9861 44863 9919 44869
rect 9861 44860 9873 44863
rect 9732 44832 9873 44860
rect 9732 44820 9738 44832
rect 9861 44829 9873 44832
rect 9907 44829 9919 44863
rect 9861 44823 9919 44829
rect 2685 44727 2743 44733
rect 2685 44693 2697 44727
rect 2731 44724 2743 44727
rect 2774 44724 2780 44736
rect 2731 44696 2780 44724
rect 2731 44693 2743 44696
rect 2685 44687 2743 44693
rect 2774 44684 2780 44696
rect 2832 44684 2838 44736
rect 10042 44724 10048 44736
rect 10003 44696 10048 44724
rect 10042 44684 10048 44696
rect 10100 44684 10106 44736
rect 1104 44634 10856 44656
rect 1104 44582 4213 44634
rect 4265 44582 4277 44634
rect 4329 44582 4341 44634
rect 4393 44582 4405 44634
rect 4457 44582 4469 44634
rect 4521 44582 7477 44634
rect 7529 44582 7541 44634
rect 7593 44582 7605 44634
rect 7657 44582 7669 44634
rect 7721 44582 7733 44634
rect 7785 44582 10856 44634
rect 1104 44560 10856 44582
rect 1486 44520 1492 44532
rect 1447 44492 1492 44520
rect 1486 44480 1492 44492
rect 1544 44480 1550 44532
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44384 1731 44387
rect 1762 44384 1768 44396
rect 1719 44356 1768 44384
rect 1719 44353 1731 44356
rect 1673 44347 1731 44353
rect 1762 44344 1768 44356
rect 1820 44344 1826 44396
rect 2133 44387 2191 44393
rect 2133 44353 2145 44387
rect 2179 44384 2191 44387
rect 2406 44384 2412 44396
rect 2179 44356 2412 44384
rect 2179 44353 2191 44356
rect 2133 44347 2191 44353
rect 2406 44344 2412 44356
rect 2464 44344 2470 44396
rect 3142 44384 3148 44396
rect 3103 44356 3148 44384
rect 3142 44344 3148 44356
rect 3200 44344 3206 44396
rect 3605 44387 3663 44393
rect 3605 44353 3617 44387
rect 3651 44353 3663 44387
rect 3605 44347 3663 44353
rect 3789 44387 3847 44393
rect 3789 44353 3801 44387
rect 3835 44384 3847 44387
rect 4154 44384 4160 44396
rect 3835 44356 4160 44384
rect 3835 44353 3847 44356
rect 3789 44347 3847 44353
rect 201 44319 259 44325
rect 201 44285 213 44319
rect 247 44316 259 44319
rect 3620 44316 3648 44347
rect 4154 44344 4160 44356
rect 4212 44344 4218 44396
rect 9766 44344 9772 44396
rect 9824 44384 9830 44396
rect 9861 44387 9919 44393
rect 9861 44384 9873 44387
rect 9824 44356 9873 44384
rect 9824 44344 9830 44356
rect 9861 44353 9873 44356
rect 9907 44353 9919 44387
rect 9861 44347 9919 44353
rect 247 44288 3648 44316
rect 3697 44319 3755 44325
rect 247 44285 259 44288
rect 201 44279 259 44285
rect 2148 44260 2176 44288
rect 3697 44285 3709 44319
rect 3743 44316 3755 44319
rect 9674 44316 9680 44328
rect 3743 44288 9680 44316
rect 3743 44285 3755 44288
rect 3697 44279 3755 44285
rect 9674 44276 9680 44288
rect 9732 44276 9738 44328
rect 2130 44208 2136 44260
rect 2188 44208 2194 44260
rect 2406 44208 2412 44260
rect 2464 44248 2470 44260
rect 5534 44248 5540 44260
rect 2464 44220 5540 44248
rect 2464 44208 2470 44220
rect 5534 44208 5540 44220
rect 5592 44208 5598 44260
rect 2314 44180 2320 44192
rect 2275 44152 2320 44180
rect 2314 44140 2320 44152
rect 2372 44140 2378 44192
rect 2958 44180 2964 44192
rect 2919 44152 2964 44180
rect 2958 44140 2964 44152
rect 3016 44140 3022 44192
rect 3234 44140 3240 44192
rect 3292 44180 3298 44192
rect 3786 44180 3792 44192
rect 3292 44152 3792 44180
rect 3292 44140 3298 44152
rect 3786 44140 3792 44152
rect 3844 44140 3850 44192
rect 10042 44180 10048 44192
rect 10003 44152 10048 44180
rect 10042 44140 10048 44152
rect 10100 44140 10106 44192
rect 1104 44090 10856 44112
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5845 44090
rect 5897 44038 5909 44090
rect 5961 44038 5973 44090
rect 6025 44038 6037 44090
rect 6089 44038 6101 44090
rect 6153 44038 9109 44090
rect 9161 44038 9173 44090
rect 9225 44038 9237 44090
rect 9289 44038 9301 44090
rect 9353 44038 9365 44090
rect 9417 44038 10856 44090
rect 1104 44016 10856 44038
rect 566 43936 572 43988
rect 624 43976 630 43988
rect 1210 43976 1216 43988
rect 624 43948 1216 43976
rect 624 43936 630 43948
rect 1210 43936 1216 43948
rect 1268 43936 1274 43988
rect 5534 43936 5540 43988
rect 5592 43976 5598 43988
rect 6178 43976 6184 43988
rect 5592 43948 6184 43976
rect 5592 43936 5598 43948
rect 6178 43936 6184 43948
rect 6236 43936 6242 43988
rect 753 43843 811 43849
rect 753 43809 765 43843
rect 799 43840 811 43843
rect 1489 43843 1547 43849
rect 1489 43840 1501 43843
rect 799 43812 1501 43840
rect 799 43809 811 43812
rect 753 43803 811 43809
rect 1489 43809 1501 43812
rect 1535 43809 1547 43843
rect 2130 43840 2136 43852
rect 1489 43803 1547 43809
rect 1596 43812 2136 43840
rect 1596 43781 1624 43812
rect 2130 43800 2136 43812
rect 2188 43840 2194 43852
rect 2498 43840 2504 43852
rect 2188 43812 2504 43840
rect 2188 43800 2194 43812
rect 2498 43800 2504 43812
rect 2556 43800 2562 43852
rect 6178 43800 6184 43852
rect 6236 43840 6242 43852
rect 6730 43840 6736 43852
rect 6236 43812 6736 43840
rect 6236 43800 6242 43812
rect 6730 43800 6736 43812
rect 6788 43800 6794 43852
rect 1581 43775 1639 43781
rect 1581 43741 1593 43775
rect 1627 43741 1639 43775
rect 1581 43735 1639 43741
rect 1670 43732 1676 43784
rect 1728 43772 1734 43784
rect 1765 43775 1823 43781
rect 1765 43772 1777 43775
rect 1728 43744 1777 43772
rect 1728 43732 1734 43744
rect 1765 43741 1777 43744
rect 1811 43741 1823 43775
rect 1765 43735 1823 43741
rect 1854 43732 1860 43784
rect 1912 43772 1918 43784
rect 2593 43775 2651 43781
rect 2593 43772 2605 43775
rect 1912 43744 2605 43772
rect 1912 43732 1918 43744
rect 2593 43741 2605 43744
rect 2639 43741 2651 43775
rect 3053 43775 3111 43781
rect 3053 43772 3065 43775
rect 2593 43735 2651 43741
rect 2746 43744 3065 43772
rect 566 43664 572 43716
rect 624 43704 630 43716
rect 2746 43704 2774 43744
rect 3053 43741 3065 43744
rect 3099 43741 3111 43775
rect 3053 43735 3111 43741
rect 3237 43775 3295 43781
rect 3237 43741 3249 43775
rect 3283 43772 3295 43775
rect 3602 43772 3608 43784
rect 3283 43744 3608 43772
rect 3283 43741 3295 43744
rect 3237 43735 3295 43741
rect 3602 43732 3608 43744
rect 3660 43772 3666 43784
rect 4154 43772 4160 43784
rect 3660 43744 4160 43772
rect 3660 43732 3666 43744
rect 4154 43732 4160 43744
rect 4212 43732 4218 43784
rect 9582 43732 9588 43784
rect 9640 43772 9646 43784
rect 9861 43775 9919 43781
rect 9861 43772 9873 43775
rect 9640 43744 9873 43772
rect 9640 43732 9646 43744
rect 9861 43741 9873 43744
rect 9907 43741 9919 43775
rect 9861 43735 9919 43741
rect 624 43676 2774 43704
rect 624 43664 630 43676
rect 2958 43664 2964 43716
rect 3016 43704 3022 43716
rect 8294 43704 8300 43716
rect 3016 43676 8300 43704
rect 3016 43664 3022 43676
rect 8294 43664 8300 43676
rect 8352 43664 8358 43716
rect 2409 43639 2467 43645
rect 2409 43605 2421 43639
rect 2455 43636 2467 43639
rect 2774 43636 2780 43648
rect 2455 43608 2780 43636
rect 2455 43605 2467 43608
rect 2409 43599 2467 43605
rect 2774 43596 2780 43608
rect 2832 43596 2838 43648
rect 3145 43639 3203 43645
rect 3145 43605 3157 43639
rect 3191 43636 3203 43639
rect 9674 43636 9680 43648
rect 3191 43608 9680 43636
rect 3191 43605 3203 43608
rect 3145 43599 3203 43605
rect 9674 43596 9680 43608
rect 9732 43596 9738 43648
rect 10042 43636 10048 43648
rect 10003 43608 10048 43636
rect 10042 43596 10048 43608
rect 10100 43596 10106 43648
rect 1104 43546 10856 43568
rect 1104 43494 4213 43546
rect 4265 43494 4277 43546
rect 4329 43494 4341 43546
rect 4393 43494 4405 43546
rect 4457 43494 4469 43546
rect 4521 43494 7477 43546
rect 7529 43494 7541 43546
rect 7593 43494 7605 43546
rect 7657 43494 7669 43546
rect 7721 43494 7733 43546
rect 7785 43494 10856 43546
rect 1104 43472 10856 43494
rect 3329 43435 3387 43441
rect 3329 43401 3341 43435
rect 3375 43432 3387 43435
rect 3878 43432 3884 43444
rect 3375 43404 3884 43432
rect 3375 43401 3387 43404
rect 3329 43395 3387 43401
rect 3878 43392 3884 43404
rect 3936 43392 3942 43444
rect 4617 43435 4675 43441
rect 4617 43401 4629 43435
rect 4663 43432 4675 43435
rect 9858 43432 9864 43444
rect 4663 43404 9864 43432
rect 4663 43401 4675 43404
rect 4617 43395 4675 43401
rect 9858 43392 9864 43404
rect 9916 43392 9922 43444
rect 934 43324 940 43376
rect 992 43364 998 43376
rect 1673 43367 1731 43373
rect 1673 43364 1685 43367
rect 992 43336 1685 43364
rect 992 43324 998 43336
rect 1673 43333 1685 43336
rect 1719 43333 1731 43367
rect 2130 43364 2136 43376
rect 1673 43327 1731 43333
rect 1872 43336 2136 43364
rect 1872 43305 1900 43336
rect 2130 43324 2136 43336
rect 2188 43324 2194 43376
rect 2958 43364 2964 43376
rect 2746 43336 2964 43364
rect 1857 43299 1915 43305
rect 1857 43265 1869 43299
rect 1903 43265 1915 43299
rect 1857 43259 1915 43265
rect 1949 43299 2007 43305
rect 1949 43265 1961 43299
rect 1995 43265 2007 43299
rect 1949 43259 2007 43265
rect 934 43188 940 43240
rect 992 43228 998 43240
rect 1118 43228 1124 43240
rect 992 43200 1124 43228
rect 992 43188 998 43200
rect 1118 43188 1124 43200
rect 1176 43228 1182 43240
rect 1964 43228 1992 43259
rect 1176 43200 1992 43228
rect 2148 43228 2176 43324
rect 2501 43299 2559 43305
rect 2501 43265 2513 43299
rect 2547 43296 2559 43299
rect 2746 43296 2774 43336
rect 2958 43324 2964 43336
rect 3016 43324 3022 43376
rect 3050 43324 3056 43376
rect 3108 43364 3114 43376
rect 3973 43367 4031 43373
rect 3108 43336 3924 43364
rect 3108 43324 3114 43336
rect 3896 43308 3924 43336
rect 3973 43333 3985 43367
rect 4019 43364 4031 43367
rect 9766 43364 9772 43376
rect 4019 43336 9772 43364
rect 4019 43333 4031 43336
rect 3973 43327 4031 43333
rect 9766 43324 9772 43336
rect 9824 43324 9830 43376
rect 2547 43268 2774 43296
rect 3237 43299 3295 43305
rect 2547 43265 2559 43268
rect 2501 43259 2559 43265
rect 3237 43265 3249 43299
rect 3283 43265 3295 43299
rect 3237 43259 3295 43265
rect 3421 43299 3479 43305
rect 3421 43265 3433 43299
rect 3467 43265 3479 43299
rect 3421 43259 3479 43265
rect 3252 43228 3280 43259
rect 2148 43200 3280 43228
rect 1176 43188 1182 43200
rect 566 43120 572 43172
rect 624 43160 630 43172
rect 3436 43160 3464 43259
rect 3602 43256 3608 43308
rect 3660 43256 3666 43308
rect 3878 43296 3884 43308
rect 3839 43268 3884 43296
rect 3878 43256 3884 43268
rect 3936 43256 3942 43308
rect 4065 43299 4123 43305
rect 4065 43265 4077 43299
rect 4111 43296 4123 43299
rect 4154 43296 4160 43308
rect 4111 43268 4160 43296
rect 4111 43265 4123 43268
rect 4065 43259 4123 43265
rect 3620 43228 3648 43256
rect 4080 43228 4108 43259
rect 4154 43256 4160 43268
rect 4212 43256 4218 43308
rect 4525 43299 4583 43305
rect 4525 43265 4537 43299
rect 4571 43265 4583 43299
rect 4525 43259 4583 43265
rect 4709 43299 4767 43305
rect 4709 43265 4721 43299
rect 4755 43265 4767 43299
rect 4709 43259 4767 43265
rect 3620 43200 4108 43228
rect 624 43132 3464 43160
rect 624 43120 630 43132
rect 3602 43120 3608 43172
rect 3660 43160 3666 43172
rect 4540 43160 4568 43259
rect 3660 43132 4568 43160
rect 3660 43120 3666 43132
rect 2685 43095 2743 43101
rect 2685 43061 2697 43095
rect 2731 43092 2743 43095
rect 2958 43092 2964 43104
rect 2731 43064 2964 43092
rect 2731 43061 2743 43064
rect 2685 43055 2743 43061
rect 2958 43052 2964 43064
rect 3016 43052 3022 43104
rect 4154 43052 4160 43104
rect 4212 43092 4218 43104
rect 4724 43092 4752 43259
rect 4212 43064 4752 43092
rect 4212 43052 4218 43064
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5845 43002
rect 5897 42950 5909 43002
rect 5961 42950 5973 43002
rect 6025 42950 6037 43002
rect 6089 42950 6101 43002
rect 6153 42950 9109 43002
rect 9161 42950 9173 43002
rect 9225 42950 9237 43002
rect 9289 42950 9301 43002
rect 9353 42950 9365 43002
rect 9417 42950 10856 43002
rect 1104 42928 10856 42950
rect 661 42891 719 42897
rect 661 42857 673 42891
rect 707 42888 719 42891
rect 1581 42891 1639 42897
rect 1581 42888 1593 42891
rect 707 42860 1593 42888
rect 707 42857 719 42860
rect 661 42851 719 42857
rect 1581 42857 1593 42860
rect 1627 42857 1639 42891
rect 4154 42888 4160 42900
rect 1581 42851 1639 42857
rect 2884 42860 4160 42888
rect 2884 42832 2912 42860
rect 2866 42780 2872 42832
rect 2924 42780 2930 42832
rect 1397 42687 1455 42693
rect 1397 42653 1409 42687
rect 1443 42653 1455 42687
rect 1397 42647 1455 42653
rect 1581 42687 1639 42693
rect 1581 42653 1593 42687
rect 1627 42684 1639 42687
rect 2130 42684 2136 42696
rect 1627 42656 2136 42684
rect 1627 42653 1639 42656
rect 1581 42647 1639 42653
rect 1412 42616 1440 42647
rect 2130 42644 2136 42656
rect 2188 42644 2194 42696
rect 2409 42687 2467 42693
rect 2409 42653 2421 42687
rect 2455 42653 2467 42687
rect 2409 42647 2467 42653
rect 2869 42687 2927 42693
rect 2869 42653 2881 42687
rect 2915 42684 2927 42687
rect 3694 42684 3700 42696
rect 2915 42656 3700 42684
rect 2915 42653 2927 42656
rect 2869 42647 2927 42653
rect 1670 42616 1676 42628
rect 1412 42588 1676 42616
rect 1670 42576 1676 42588
rect 1728 42576 1734 42628
rect 2424 42616 2452 42647
rect 3694 42644 3700 42656
rect 3752 42644 3758 42696
rect 3988 42693 4016 42860
rect 4154 42848 4160 42860
rect 4212 42848 4218 42900
rect 9674 42780 9680 42832
rect 9732 42820 9738 42832
rect 9732 42792 9904 42820
rect 9732 42780 9738 42792
rect 9876 42693 9904 42792
rect 3789 42687 3847 42693
rect 3789 42653 3801 42687
rect 3835 42653 3847 42687
rect 3789 42647 3847 42653
rect 3973 42687 4031 42693
rect 3973 42653 3985 42687
rect 4019 42653 4031 42687
rect 3973 42647 4031 42653
rect 9861 42687 9919 42693
rect 9861 42653 9873 42687
rect 9907 42653 9919 42687
rect 9861 42647 9919 42653
rect 2498 42616 2504 42628
rect 2424 42588 2504 42616
rect 2498 42576 2504 42588
rect 2556 42616 2562 42628
rect 3804 42616 3832 42647
rect 2556 42588 3832 42616
rect 3881 42619 3939 42625
rect 2556 42576 2562 42588
rect 3881 42585 3893 42619
rect 3927 42616 3939 42619
rect 10965 42619 11023 42625
rect 10965 42616 10977 42619
rect 3927 42588 10977 42616
rect 3927 42585 3939 42588
rect 3881 42579 3939 42585
rect 10965 42585 10977 42588
rect 11011 42585 11023 42619
rect 10965 42579 11023 42585
rect 842 42508 848 42560
rect 900 42548 906 42560
rect 2133 42551 2191 42557
rect 2133 42548 2145 42551
rect 900 42520 2145 42548
rect 900 42508 906 42520
rect 2133 42517 2145 42520
rect 2179 42517 2191 42551
rect 3050 42548 3056 42560
rect 3011 42520 3056 42548
rect 2133 42511 2191 42517
rect 3050 42508 3056 42520
rect 3108 42508 3114 42560
rect 10042 42548 10048 42560
rect 10003 42520 10048 42548
rect 10042 42508 10048 42520
rect 10100 42508 10106 42560
rect 1104 42458 10856 42480
rect 1104 42406 4213 42458
rect 4265 42406 4277 42458
rect 4329 42406 4341 42458
rect 4393 42406 4405 42458
rect 4457 42406 4469 42458
rect 4521 42406 7477 42458
rect 7529 42406 7541 42458
rect 7593 42406 7605 42458
rect 7657 42406 7669 42458
rect 7721 42406 7733 42458
rect 7785 42406 10856 42458
rect 1104 42384 10856 42406
rect 3237 42347 3295 42353
rect 3237 42313 3249 42347
rect 3283 42344 3295 42347
rect 9582 42344 9588 42356
rect 3283 42316 9588 42344
rect 3283 42313 3295 42316
rect 3237 42307 3295 42313
rect 9582 42304 9588 42316
rect 9640 42304 9646 42356
rect 1688 42248 2912 42276
rect 1688 42217 1716 42248
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42177 1731 42211
rect 2406 42208 2412 42220
rect 2367 42180 2412 42208
rect 1673 42171 1731 42177
rect 2406 42168 2412 42180
rect 2464 42168 2470 42220
rect 2884 42140 2912 42248
rect 2958 42236 2964 42288
rect 3016 42276 3022 42288
rect 3016 42248 3372 42276
rect 3016 42236 3022 42248
rect 3344 42217 3372 42248
rect 3053 42211 3111 42217
rect 3053 42177 3065 42211
rect 3099 42208 3111 42211
rect 3145 42211 3203 42217
rect 3145 42208 3157 42211
rect 3099 42180 3157 42208
rect 3099 42177 3111 42180
rect 3053 42171 3111 42177
rect 3145 42177 3157 42180
rect 3191 42177 3203 42211
rect 3145 42171 3203 42177
rect 3329 42211 3387 42217
rect 3329 42177 3341 42211
rect 3375 42177 3387 42211
rect 9858 42208 9864 42220
rect 9819 42180 9864 42208
rect 3329 42171 3387 42177
rect 9858 42168 9864 42180
rect 9916 42168 9922 42220
rect 11333 42143 11391 42149
rect 11333 42140 11345 42143
rect 2884 42112 11345 42140
rect 11333 42109 11345 42112
rect 11379 42109 11391 42143
rect 11333 42103 11391 42109
rect 1670 42032 1676 42084
rect 1728 42072 1734 42084
rect 1728 42044 2360 42072
rect 1728 42032 1734 42044
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 2222 42004 2228 42016
rect 2183 41976 2228 42004
rect 2222 41964 2228 41976
rect 2280 41964 2286 42016
rect 2332 42004 2360 42044
rect 3053 42007 3111 42013
rect 3053 42004 3065 42007
rect 2332 41976 3065 42004
rect 3053 41973 3065 41976
rect 3099 41973 3111 42007
rect 10042 42004 10048 42016
rect 10003 41976 10048 42004
rect 3053 41967 3111 41973
rect 10042 41964 10048 41976
rect 10100 41964 10106 42016
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5845 41914
rect 5897 41862 5909 41914
rect 5961 41862 5973 41914
rect 6025 41862 6037 41914
rect 6089 41862 6101 41914
rect 6153 41862 9109 41914
rect 9161 41862 9173 41914
rect 9225 41862 9237 41914
rect 9289 41862 9301 41914
rect 9353 41862 9365 41914
rect 9417 41862 10856 41914
rect 1104 41840 10856 41862
rect 2961 41803 3019 41809
rect 2961 41769 2973 41803
rect 3007 41800 3019 41803
rect 9858 41800 9864 41812
rect 3007 41772 9864 41800
rect 3007 41769 3019 41772
rect 2961 41763 3019 41769
rect 9858 41760 9864 41772
rect 9916 41760 9922 41812
rect 1854 41692 1860 41744
rect 1912 41732 1918 41744
rect 3786 41732 3792 41744
rect 1912 41704 3792 41732
rect 1912 41692 1918 41704
rect 3786 41692 3792 41704
rect 3844 41692 3850 41744
rect 198 41624 204 41676
rect 256 41664 262 41676
rect 1949 41667 2007 41673
rect 1949 41664 1961 41667
rect 256 41636 1961 41664
rect 256 41624 262 41636
rect 1949 41633 1961 41636
rect 1995 41633 2007 41667
rect 1949 41627 2007 41633
rect 2222 41624 2228 41676
rect 2280 41664 2286 41676
rect 2280 41636 2464 41664
rect 2280 41624 2286 41636
rect 937 41599 995 41605
rect 937 41565 949 41599
rect 983 41596 995 41599
rect 1762 41596 1768 41608
rect 983 41568 1768 41596
rect 983 41565 995 41568
rect 937 41559 995 41565
rect 1762 41556 1768 41568
rect 1820 41556 1826 41608
rect 1854 41556 1860 41608
rect 1912 41596 1918 41608
rect 2130 41596 2136 41608
rect 1912 41568 1992 41596
rect 2091 41568 2136 41596
rect 1912 41556 1918 41568
rect 198 41528 204 41540
rect 159 41500 204 41528
rect 198 41488 204 41500
rect 256 41488 262 41540
rect 1029 41531 1087 41537
rect 1029 41497 1041 41531
rect 1075 41528 1087 41531
rect 1964 41528 1992 41568
rect 2130 41556 2136 41568
rect 2188 41556 2194 41608
rect 2317 41599 2375 41605
rect 2317 41565 2329 41599
rect 2363 41565 2375 41599
rect 2436 41596 2464 41636
rect 2682 41624 2688 41676
rect 2740 41664 2746 41676
rect 7006 41664 7012 41676
rect 2740 41636 7012 41664
rect 2740 41624 2746 41636
rect 7006 41624 7012 41636
rect 7064 41624 7070 41676
rect 2777 41599 2835 41605
rect 2777 41596 2789 41599
rect 2436 41568 2789 41596
rect 2317 41559 2375 41565
rect 2777 41565 2789 41568
rect 2823 41565 2835 41599
rect 2958 41596 2964 41608
rect 2919 41568 2964 41596
rect 2777 41559 2835 41565
rect 2332 41528 2360 41559
rect 2958 41556 2964 41568
rect 3016 41556 3022 41608
rect 3602 41528 3608 41540
rect 1075 41500 1900 41528
rect 1964 41500 3608 41528
rect 1075 41497 1087 41500
rect 1029 41491 1087 41497
rect 1210 41420 1216 41472
rect 1268 41460 1274 41472
rect 1762 41460 1768 41472
rect 1268 41432 1768 41460
rect 1268 41420 1274 41432
rect 1762 41420 1768 41432
rect 1820 41420 1826 41472
rect 1872 41460 1900 41500
rect 3602 41488 3608 41500
rect 3660 41488 3666 41540
rect 2406 41460 2412 41472
rect 1872 41432 2412 41460
rect 2406 41420 2412 41432
rect 2464 41420 2470 41472
rect 3418 41420 3424 41472
rect 3476 41460 3482 41472
rect 5718 41460 5724 41472
rect 3476 41432 5724 41460
rect 3476 41420 3482 41432
rect 5718 41420 5724 41432
rect 5776 41420 5782 41472
rect 1104 41370 10856 41392
rect 1104 41318 4213 41370
rect 4265 41318 4277 41370
rect 4329 41318 4341 41370
rect 4393 41318 4405 41370
rect 4457 41318 4469 41370
rect 4521 41318 7477 41370
rect 7529 41318 7541 41370
rect 7593 41318 7605 41370
rect 7657 41318 7669 41370
rect 7721 41318 7733 41370
rect 7785 41318 10856 41370
rect 1104 41296 10856 41318
rect 3326 41216 3332 41268
rect 3384 41256 3390 41268
rect 3970 41256 3976 41268
rect 3384 41228 3976 41256
rect 3384 41216 3390 41228
rect 3970 41216 3976 41228
rect 4028 41216 4034 41268
rect 8386 41188 8392 41200
rect 1688 41160 8392 41188
rect 1688 41129 1716 41160
rect 8386 41148 8392 41160
rect 8444 41148 8450 41200
rect 1673 41123 1731 41129
rect 1673 41089 1685 41123
rect 1719 41089 1731 41123
rect 1673 41083 1731 41089
rect 2409 41123 2467 41129
rect 2409 41089 2421 41123
rect 2455 41120 2467 41123
rect 2682 41120 2688 41132
rect 2455 41092 2688 41120
rect 2455 41089 2467 41092
rect 2409 41083 2467 41089
rect 2682 41080 2688 41092
rect 2740 41080 2746 41132
rect 2869 41123 2927 41129
rect 2869 41089 2881 41123
rect 2915 41120 2927 41123
rect 4062 41120 4068 41132
rect 2915 41092 4068 41120
rect 2915 41089 2927 41092
rect 2869 41083 2927 41089
rect 4062 41080 4068 41092
rect 4120 41080 4126 41132
rect 9674 41080 9680 41132
rect 9732 41120 9738 41132
rect 9861 41123 9919 41129
rect 9861 41120 9873 41123
rect 9732 41092 9873 41120
rect 9732 41080 9738 41092
rect 9861 41089 9873 41092
rect 9907 41089 9919 41123
rect 9861 41083 9919 41089
rect 2038 41012 2044 41064
rect 2096 41052 2102 41064
rect 2222 41052 2228 41064
rect 2096 41024 2228 41052
rect 2096 41012 2102 41024
rect 2222 41012 2228 41024
rect 2280 41012 2286 41064
rect 3050 40984 3056 40996
rect 3011 40956 3056 40984
rect 3050 40944 3056 40956
rect 3108 40944 3114 40996
rect 10042 40984 10048 40996
rect 10003 40956 10048 40984
rect 10042 40944 10048 40956
rect 10100 40944 10106 40996
rect 1210 40876 1216 40928
rect 1268 40916 1274 40928
rect 1489 40919 1547 40925
rect 1489 40916 1501 40919
rect 1268 40888 1501 40916
rect 1268 40876 1274 40888
rect 1489 40885 1501 40888
rect 1535 40885 1547 40919
rect 2222 40916 2228 40928
rect 2183 40888 2228 40916
rect 1489 40879 1547 40885
rect 2222 40876 2228 40888
rect 2280 40876 2286 40928
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5845 40826
rect 5897 40774 5909 40826
rect 5961 40774 5973 40826
rect 6025 40774 6037 40826
rect 6089 40774 6101 40826
rect 6153 40774 9109 40826
rect 9161 40774 9173 40826
rect 9225 40774 9237 40826
rect 9289 40774 9301 40826
rect 9353 40774 9365 40826
rect 9417 40774 10856 40826
rect 1104 40752 10856 40774
rect 658 40672 664 40724
rect 716 40712 722 40724
rect 2133 40715 2191 40721
rect 2133 40712 2145 40715
rect 716 40684 2145 40712
rect 716 40672 722 40684
rect 2133 40681 2145 40684
rect 2179 40681 2191 40715
rect 2133 40675 2191 40681
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 1762 40508 1768 40520
rect 1719 40480 1768 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 1762 40468 1768 40480
rect 1820 40468 1826 40520
rect 2133 40511 2191 40517
rect 2133 40477 2145 40511
rect 2179 40477 2191 40511
rect 2133 40471 2191 40477
rect 2317 40511 2375 40517
rect 2317 40477 2329 40511
rect 2363 40508 2375 40511
rect 2866 40508 2872 40520
rect 2363 40480 2872 40508
rect 2363 40477 2375 40480
rect 2317 40471 2375 40477
rect 2148 40440 2176 40471
rect 2866 40468 2872 40480
rect 2924 40468 2930 40520
rect 9858 40508 9864 40520
rect 9819 40480 9864 40508
rect 9858 40468 9864 40480
rect 9916 40468 9922 40520
rect 2590 40440 2596 40452
rect 2148 40412 2596 40440
rect 2590 40400 2596 40412
rect 2648 40400 2654 40452
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 10042 40372 10048 40384
rect 10003 40344 10048 40372
rect 10042 40332 10048 40344
rect 10100 40332 10106 40384
rect 1104 40282 10856 40304
rect 1104 40230 4213 40282
rect 4265 40230 4277 40282
rect 4329 40230 4341 40282
rect 4393 40230 4405 40282
rect 4457 40230 4469 40282
rect 4521 40230 7477 40282
rect 7529 40230 7541 40282
rect 7593 40230 7605 40282
rect 7657 40230 7669 40282
rect 7721 40230 7733 40282
rect 7785 40230 10856 40282
rect 1104 40208 10856 40230
rect 1854 40128 1860 40180
rect 1912 40168 1918 40180
rect 2590 40168 2596 40180
rect 1912 40140 2596 40168
rect 1912 40128 1918 40140
rect 2590 40128 2596 40140
rect 2648 40128 2654 40180
rect 2225 40103 2283 40109
rect 2225 40069 2237 40103
rect 2271 40100 2283 40103
rect 4798 40100 4804 40112
rect 2271 40072 4804 40100
rect 2271 40069 2283 40072
rect 2225 40063 2283 40069
rect 4798 40060 4804 40072
rect 4856 40060 4862 40112
rect 845 40035 903 40041
rect 845 40001 857 40035
rect 891 40032 903 40035
rect 1673 40035 1731 40041
rect 1673 40032 1685 40035
rect 891 40004 1685 40032
rect 891 40001 903 40004
rect 845 39995 903 40001
rect 1673 40001 1685 40004
rect 1719 40001 1731 40035
rect 1673 39995 1731 40001
rect 1854 39992 1860 40044
rect 1912 40032 1918 40044
rect 2133 40035 2191 40041
rect 2133 40032 2145 40035
rect 1912 40004 2145 40032
rect 1912 39992 1918 40004
rect 2133 40001 2145 40004
rect 2179 40001 2191 40035
rect 2133 39995 2191 40001
rect 2314 39992 2320 40044
rect 2372 40032 2378 40044
rect 2866 40032 2872 40044
rect 2372 40004 2465 40032
rect 2827 40004 2872 40032
rect 2372 39992 2378 40004
rect 2866 39992 2872 40004
rect 2924 39992 2930 40044
rect 3050 40032 3056 40044
rect 3011 40004 3056 40032
rect 3050 39992 3056 40004
rect 3108 39992 3114 40044
rect 9766 39992 9772 40044
rect 9824 40032 9830 40044
rect 9861 40035 9919 40041
rect 9861 40032 9873 40035
rect 9824 40004 9873 40032
rect 9824 39992 9830 40004
rect 9861 40001 9873 40004
rect 9907 40001 9919 40035
rect 9861 39995 9919 40001
rect 2332 39964 2360 39992
rect 2056 39936 2360 39964
rect 1210 39788 1216 39840
rect 1268 39828 1274 39840
rect 1489 39831 1547 39837
rect 1489 39828 1501 39831
rect 1268 39800 1501 39828
rect 1268 39788 1274 39800
rect 1489 39797 1501 39800
rect 1535 39797 1547 39831
rect 2056 39828 2084 39936
rect 3053 39899 3111 39905
rect 3053 39865 3065 39899
rect 3099 39896 3111 39899
rect 9674 39896 9680 39908
rect 3099 39868 9680 39896
rect 3099 39865 3111 39868
rect 3053 39859 3111 39865
rect 9674 39856 9680 39868
rect 9732 39856 9738 39908
rect 2222 39828 2228 39840
rect 2056 39800 2228 39828
rect 1489 39791 1547 39797
rect 2222 39788 2228 39800
rect 2280 39788 2286 39840
rect 10042 39828 10048 39840
rect 10003 39800 10048 39828
rect 10042 39788 10048 39800
rect 10100 39788 10106 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5845 39738
rect 5897 39686 5909 39738
rect 5961 39686 5973 39738
rect 6025 39686 6037 39738
rect 6089 39686 6101 39738
rect 6153 39686 9109 39738
rect 9161 39686 9173 39738
rect 9225 39686 9237 39738
rect 9289 39686 9301 39738
rect 9353 39686 9365 39738
rect 9417 39686 10856 39738
rect 1104 39664 10856 39686
rect 14 39448 20 39500
rect 72 39488 78 39500
rect 1581 39491 1639 39497
rect 1581 39488 1593 39491
rect 72 39460 1593 39488
rect 72 39448 78 39460
rect 1581 39457 1593 39460
rect 1627 39457 1639 39491
rect 1581 39451 1639 39457
rect 1486 39380 1492 39432
rect 1544 39420 1550 39432
rect 1673 39423 1731 39429
rect 1673 39420 1685 39423
rect 1544 39392 1685 39420
rect 1544 39380 1550 39392
rect 1673 39389 1685 39392
rect 1719 39420 1731 39423
rect 1854 39420 1860 39432
rect 1719 39392 1860 39420
rect 1719 39389 1731 39392
rect 1673 39383 1731 39389
rect 1854 39380 1860 39392
rect 1912 39380 1918 39432
rect 1949 39423 2007 39429
rect 1949 39389 1961 39423
rect 1995 39389 2007 39423
rect 1949 39383 2007 39389
rect 2409 39423 2467 39429
rect 2409 39389 2421 39423
rect 2455 39420 2467 39423
rect 3418 39420 3424 39432
rect 2455 39392 3424 39420
rect 2455 39389 2467 39392
rect 2409 39383 2467 39389
rect 1964 39352 1992 39383
rect 3418 39380 3424 39392
rect 3476 39380 3482 39432
rect 2866 39352 2872 39364
rect 1964 39324 2872 39352
rect 2866 39312 2872 39324
rect 2924 39312 2930 39364
rect 2593 39287 2651 39293
rect 2593 39253 2605 39287
rect 2639 39284 2651 39287
rect 2774 39284 2780 39296
rect 2639 39256 2780 39284
rect 2639 39253 2651 39256
rect 2593 39247 2651 39253
rect 2774 39244 2780 39256
rect 2832 39244 2838 39296
rect 1104 39194 10856 39216
rect 1104 39142 4213 39194
rect 4265 39142 4277 39194
rect 4329 39142 4341 39194
rect 4393 39142 4405 39194
rect 4457 39142 4469 39194
rect 4521 39142 7477 39194
rect 7529 39142 7541 39194
rect 7593 39142 7605 39194
rect 7657 39142 7669 39194
rect 7721 39142 7733 39194
rect 7785 39142 10856 39194
rect 1104 39120 10856 39142
rect 1949 39083 2007 39089
rect 1949 39049 1961 39083
rect 1995 39080 2007 39083
rect 3510 39080 3516 39092
rect 1995 39052 3516 39080
rect 1995 39049 2007 39052
rect 1949 39043 2007 39049
rect 3510 39040 3516 39052
rect 3568 39040 3574 39092
rect 4065 39083 4123 39089
rect 4065 39049 4077 39083
rect 4111 39080 4123 39083
rect 9858 39080 9864 39092
rect 4111 39052 9864 39080
rect 4111 39049 4123 39052
rect 4065 39043 4123 39049
rect 9858 39040 9864 39052
rect 9916 39040 9922 39092
rect 3602 39012 3608 39024
rect 2792 38984 3608 39012
rect 1854 38944 1860 38956
rect 1815 38916 1860 38944
rect 1854 38904 1860 38916
rect 1912 38904 1918 38956
rect 2792 38953 2820 38984
rect 3602 38972 3608 38984
rect 3660 38972 3666 39024
rect 2777 38947 2835 38953
rect 2777 38913 2789 38947
rect 2823 38913 2835 38947
rect 3234 38944 3240 38956
rect 3195 38916 3240 38944
rect 2777 38907 2835 38913
rect 3234 38904 3240 38916
rect 3292 38904 3298 38956
rect 3973 38947 4031 38953
rect 3973 38913 3985 38947
rect 4019 38913 4031 38947
rect 3973 38907 4031 38913
rect 2958 38836 2964 38888
rect 3016 38876 3022 38888
rect 3510 38876 3516 38888
rect 3016 38848 3516 38876
rect 3016 38836 3022 38848
rect 3510 38836 3516 38848
rect 3568 38836 3574 38888
rect 2866 38768 2872 38820
rect 2924 38808 2930 38820
rect 3234 38808 3240 38820
rect 2924 38780 3240 38808
rect 2924 38768 2930 38780
rect 3234 38768 3240 38780
rect 3292 38808 3298 38820
rect 3988 38808 4016 38907
rect 4062 38904 4068 38956
rect 4120 38944 4126 38956
rect 4157 38947 4215 38953
rect 4157 38944 4169 38947
rect 4120 38916 4169 38944
rect 4120 38904 4126 38916
rect 4157 38913 4169 38916
rect 4203 38913 4215 38947
rect 9858 38944 9864 38956
rect 9819 38916 9864 38944
rect 4157 38907 4215 38913
rect 9858 38904 9864 38916
rect 9916 38904 9922 38956
rect 3292 38780 4016 38808
rect 3292 38768 3298 38780
rect 2593 38743 2651 38749
rect 2593 38709 2605 38743
rect 2639 38740 2651 38743
rect 2958 38740 2964 38752
rect 2639 38712 2964 38740
rect 2639 38709 2651 38712
rect 2593 38703 2651 38709
rect 2958 38700 2964 38712
rect 3016 38700 3022 38752
rect 3418 38740 3424 38752
rect 3379 38712 3424 38740
rect 3418 38700 3424 38712
rect 3476 38700 3482 38752
rect 3694 38700 3700 38752
rect 3752 38740 3758 38752
rect 6362 38740 6368 38752
rect 3752 38712 6368 38740
rect 3752 38700 3758 38712
rect 6362 38700 6368 38712
rect 6420 38700 6426 38752
rect 10042 38740 10048 38752
rect 10003 38712 10048 38740
rect 10042 38700 10048 38712
rect 10100 38700 10106 38752
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5845 38650
rect 5897 38598 5909 38650
rect 5961 38598 5973 38650
rect 6025 38598 6037 38650
rect 6089 38598 6101 38650
rect 6153 38598 9109 38650
rect 9161 38598 9173 38650
rect 9225 38598 9237 38650
rect 9289 38598 9301 38650
rect 9353 38598 9365 38650
rect 9417 38598 10856 38650
rect 1104 38576 10856 38598
rect 1118 38496 1124 38548
rect 1176 38536 1182 38548
rect 3145 38539 3203 38545
rect 1176 38508 2452 38536
rect 1176 38496 1182 38508
rect 1486 38360 1492 38412
rect 1544 38400 1550 38412
rect 2130 38400 2136 38412
rect 1544 38372 1808 38400
rect 2091 38372 2136 38400
rect 1544 38360 1550 38372
rect 1673 38335 1731 38341
rect 1673 38332 1685 38335
rect 1596 38304 1685 38332
rect 1486 38196 1492 38208
rect 1447 38168 1492 38196
rect 1486 38156 1492 38168
rect 1544 38156 1550 38208
rect 1596 38196 1624 38304
rect 1673 38301 1685 38304
rect 1719 38301 1731 38335
rect 1780 38332 1808 38372
rect 2130 38360 2136 38372
rect 2188 38360 2194 38412
rect 2424 38341 2452 38508
rect 3145 38505 3157 38539
rect 3191 38536 3203 38539
rect 9766 38536 9772 38548
rect 3191 38508 9772 38536
rect 3191 38505 3203 38508
rect 3145 38499 3203 38505
rect 9766 38496 9772 38508
rect 9824 38496 9830 38548
rect 11333 38471 11391 38477
rect 11333 38468 11345 38471
rect 2884 38440 11345 38468
rect 2225 38335 2283 38341
rect 2225 38332 2237 38335
rect 1780 38304 2237 38332
rect 1673 38295 1731 38301
rect 2225 38301 2237 38304
rect 2271 38301 2283 38335
rect 2225 38295 2283 38301
rect 2409 38335 2467 38341
rect 2409 38301 2421 38335
rect 2455 38301 2467 38335
rect 2409 38295 2467 38301
rect 2130 38224 2136 38276
rect 2188 38264 2194 38276
rect 2240 38264 2268 38295
rect 2188 38236 2268 38264
rect 2188 38224 2194 38236
rect 2884 38196 2912 38440
rect 11333 38437 11345 38440
rect 11379 38437 11391 38471
rect 11333 38431 11391 38437
rect 3881 38403 3939 38409
rect 3881 38369 3893 38403
rect 3927 38400 3939 38403
rect 3927 38372 9904 38400
rect 3927 38369 3939 38372
rect 3881 38363 3939 38369
rect 2961 38335 3019 38341
rect 2961 38301 2973 38335
rect 3007 38301 3019 38335
rect 2961 38295 3019 38301
rect 1596 38168 2912 38196
rect 2976 38196 3004 38295
rect 3050 38292 3056 38344
rect 3108 38332 3114 38344
rect 3145 38335 3203 38341
rect 3145 38332 3157 38335
rect 3108 38304 3157 38332
rect 3108 38292 3114 38304
rect 3145 38301 3157 38304
rect 3191 38301 3203 38335
rect 3145 38295 3203 38301
rect 3160 38264 3188 38295
rect 3602 38292 3608 38344
rect 3660 38332 3666 38344
rect 3789 38335 3847 38341
rect 3789 38332 3801 38335
rect 3660 38304 3801 38332
rect 3660 38292 3666 38304
rect 3789 38301 3801 38304
rect 3835 38301 3847 38335
rect 3789 38295 3847 38301
rect 3973 38335 4031 38341
rect 3973 38301 3985 38335
rect 4019 38332 4031 38335
rect 4062 38332 4068 38344
rect 4019 38304 4068 38332
rect 4019 38301 4031 38304
rect 3973 38295 4031 38301
rect 3988 38264 4016 38295
rect 4062 38292 4068 38304
rect 4120 38292 4126 38344
rect 9876 38341 9904 38372
rect 9861 38335 9919 38341
rect 9861 38301 9873 38335
rect 9907 38301 9919 38335
rect 9861 38295 9919 38301
rect 3160 38236 4016 38264
rect 3418 38196 3424 38208
rect 2976 38168 3424 38196
rect 3418 38156 3424 38168
rect 3476 38156 3482 38208
rect 10042 38196 10048 38208
rect 10003 38168 10048 38196
rect 10042 38156 10048 38168
rect 10100 38156 10106 38208
rect 1104 38106 10856 38128
rect 1104 38054 4213 38106
rect 4265 38054 4277 38106
rect 4329 38054 4341 38106
rect 4393 38054 4405 38106
rect 4457 38054 4469 38106
rect 4521 38054 7477 38106
rect 7529 38054 7541 38106
rect 7593 38054 7605 38106
rect 7657 38054 7669 38106
rect 7721 38054 7733 38106
rect 7785 38054 10856 38106
rect 1104 38032 10856 38054
rect 750 37952 756 38004
rect 808 37992 814 38004
rect 2225 37995 2283 38001
rect 2225 37992 2237 37995
rect 808 37964 2237 37992
rect 808 37952 814 37964
rect 2225 37961 2237 37964
rect 2271 37961 2283 37995
rect 2225 37955 2283 37961
rect 3237 37995 3295 38001
rect 3237 37961 3249 37995
rect 3283 37992 3295 37995
rect 4890 37992 4896 38004
rect 3283 37964 4896 37992
rect 3283 37961 3295 37964
rect 3237 37955 3295 37961
rect 4890 37952 4896 37964
rect 4948 37952 4954 38004
rect 11149 37927 11207 37933
rect 11149 37924 11161 37927
rect 1688 37896 11161 37924
rect 1688 37865 1716 37896
rect 11149 37893 11161 37896
rect 11195 37893 11207 37927
rect 11149 37887 11207 37893
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 2130 37816 2136 37868
rect 2188 37856 2194 37868
rect 2225 37859 2283 37865
rect 2225 37856 2237 37859
rect 2188 37828 2237 37856
rect 2188 37816 2194 37828
rect 2225 37825 2237 37828
rect 2271 37825 2283 37859
rect 2225 37819 2283 37825
rect 2501 37859 2559 37865
rect 2501 37825 2513 37859
rect 2547 37825 2559 37859
rect 2501 37819 2559 37825
rect 2516 37788 2544 37819
rect 2958 37816 2964 37868
rect 3016 37856 3022 37868
rect 3053 37859 3111 37865
rect 3053 37856 3065 37859
rect 3016 37828 3065 37856
rect 3016 37816 3022 37828
rect 3053 37825 3065 37828
rect 3099 37825 3111 37859
rect 3053 37819 3111 37825
rect 3329 37859 3387 37865
rect 3329 37825 3341 37859
rect 3375 37856 3387 37859
rect 3418 37856 3424 37868
rect 3375 37828 3424 37856
rect 3375 37825 3387 37828
rect 3329 37819 3387 37825
rect 3418 37816 3424 37828
rect 3476 37816 3482 37868
rect 3602 37788 3608 37800
rect 2516 37760 3608 37788
rect 3602 37748 3608 37760
rect 3660 37748 3666 37800
rect 1486 37652 1492 37664
rect 1447 37624 1492 37652
rect 1486 37612 1492 37624
rect 1544 37612 1550 37664
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5845 37562
rect 5897 37510 5909 37562
rect 5961 37510 5973 37562
rect 6025 37510 6037 37562
rect 6089 37510 6101 37562
rect 6153 37510 9109 37562
rect 9161 37510 9173 37562
rect 9225 37510 9237 37562
rect 9289 37510 9301 37562
rect 9353 37510 9365 37562
rect 9417 37510 10856 37562
rect 1104 37488 10856 37510
rect 2130 37380 2136 37392
rect 1688 37352 2136 37380
rect 1026 37204 1032 37256
rect 1084 37244 1090 37256
rect 1688 37253 1716 37352
rect 2130 37340 2136 37352
rect 2188 37380 2194 37392
rect 2958 37380 2964 37392
rect 2188 37352 2964 37380
rect 2188 37340 2194 37352
rect 2958 37340 2964 37352
rect 3016 37340 3022 37392
rect 9858 37340 9864 37392
rect 9916 37340 9922 37392
rect 2593 37315 2651 37321
rect 2593 37281 2605 37315
rect 2639 37312 2651 37315
rect 9876 37312 9904 37340
rect 2639 37284 9904 37312
rect 2639 37281 2651 37284
rect 2593 37275 2651 37281
rect 1489 37247 1547 37253
rect 1489 37244 1501 37247
rect 1084 37216 1501 37244
rect 1084 37204 1090 37216
rect 1489 37213 1501 37216
rect 1535 37213 1547 37247
rect 1489 37207 1547 37213
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37213 1731 37247
rect 2501 37247 2559 37253
rect 2501 37244 2513 37247
rect 1673 37207 1731 37213
rect 1780 37216 2513 37244
rect 1504 37176 1532 37207
rect 1780 37176 1808 37216
rect 2501 37213 2513 37216
rect 2547 37213 2559 37247
rect 2501 37207 2559 37213
rect 2685 37247 2743 37253
rect 2685 37213 2697 37247
rect 2731 37244 2743 37247
rect 3050 37244 3056 37256
rect 2731 37216 3056 37244
rect 2731 37213 2743 37216
rect 2685 37207 2743 37213
rect 3050 37204 3056 37216
rect 3108 37204 3114 37256
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 3292 37216 9873 37244
rect 3292 37204 3298 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 1504 37148 1808 37176
rect 1857 37179 1915 37185
rect 1857 37145 1869 37179
rect 1903 37176 1915 37179
rect 4614 37176 4620 37188
rect 1903 37148 4620 37176
rect 1903 37145 1915 37148
rect 1857 37139 1915 37145
rect 4614 37136 4620 37148
rect 4672 37136 4678 37188
rect 10042 37108 10048 37120
rect 10003 37080 10048 37108
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 1104 37018 10856 37040
rect 1104 36966 4213 37018
rect 4265 36966 4277 37018
rect 4329 36966 4341 37018
rect 4393 36966 4405 37018
rect 4457 36966 4469 37018
rect 4521 36966 7477 37018
rect 7529 36966 7541 37018
rect 7593 36966 7605 37018
rect 7657 36966 7669 37018
rect 7721 36966 7733 37018
rect 7785 36966 10856 37018
rect 1104 36944 10856 36966
rect 753 36839 811 36845
rect 753 36805 765 36839
rect 799 36836 811 36839
rect 2314 36836 2320 36848
rect 799 36808 2320 36836
rect 799 36805 811 36808
rect 753 36799 811 36805
rect 2314 36796 2320 36808
rect 2372 36796 2378 36848
rect 6914 36836 6920 36848
rect 2746 36808 6920 36836
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36737 1731 36771
rect 1673 36731 1731 36737
rect 2133 36771 2191 36777
rect 2133 36737 2145 36771
rect 2179 36768 2191 36771
rect 2746 36768 2774 36808
rect 6914 36796 6920 36808
rect 6972 36796 6978 36848
rect 11057 36839 11115 36845
rect 11057 36836 11069 36839
rect 9692 36808 11069 36836
rect 2179 36740 2774 36768
rect 2869 36771 2927 36777
rect 2179 36737 2191 36740
rect 2133 36731 2191 36737
rect 2869 36737 2881 36771
rect 2915 36768 2927 36771
rect 9692 36768 9720 36808
rect 11057 36805 11069 36808
rect 11103 36805 11115 36839
rect 11057 36799 11115 36805
rect 2915 36740 9720 36768
rect 2915 36737 2927 36740
rect 2869 36731 2927 36737
rect 566 36660 572 36712
rect 624 36700 630 36712
rect 1210 36700 1216 36712
rect 624 36672 1216 36700
rect 624 36660 630 36672
rect 1210 36660 1216 36672
rect 1268 36660 1274 36712
rect 1688 36700 1716 36731
rect 9766 36728 9772 36780
rect 9824 36768 9830 36780
rect 9861 36771 9919 36777
rect 9861 36768 9873 36771
rect 9824 36740 9873 36768
rect 9824 36728 9830 36740
rect 9861 36737 9873 36740
rect 9907 36737 9919 36771
rect 9861 36731 9919 36737
rect 8478 36700 8484 36712
rect 1688 36672 8484 36700
rect 8478 36660 8484 36672
rect 8536 36660 8542 36712
rect 3050 36632 3056 36644
rect 3011 36604 3056 36632
rect 3050 36592 3056 36604
rect 3108 36592 3114 36644
rect 198 36524 204 36576
rect 256 36564 262 36576
rect 566 36564 572 36576
rect 256 36536 572 36564
rect 256 36524 262 36536
rect 566 36524 572 36536
rect 624 36524 630 36576
rect 1486 36564 1492 36576
rect 1447 36536 1492 36564
rect 1486 36524 1492 36536
rect 1544 36524 1550 36576
rect 2314 36564 2320 36576
rect 2275 36536 2320 36564
rect 2314 36524 2320 36536
rect 2372 36524 2378 36576
rect 10042 36564 10048 36576
rect 10003 36536 10048 36564
rect 10042 36524 10048 36536
rect 10100 36524 10106 36576
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5845 36474
rect 5897 36422 5909 36474
rect 5961 36422 5973 36474
rect 6025 36422 6037 36474
rect 6089 36422 6101 36474
rect 6153 36422 9109 36474
rect 9161 36422 9173 36474
rect 9225 36422 9237 36474
rect 9289 36422 9301 36474
rect 9353 36422 9365 36474
rect 9417 36422 10856 36474
rect 1104 36400 10856 36422
rect 3234 36360 3240 36372
rect 3195 36332 3240 36360
rect 3234 36320 3240 36332
rect 3292 36320 3298 36372
rect 1857 36295 1915 36301
rect 1857 36261 1869 36295
rect 1903 36292 1915 36295
rect 4982 36292 4988 36304
rect 1903 36264 4988 36292
rect 1903 36261 1915 36264
rect 1857 36255 1915 36261
rect 4982 36252 4988 36264
rect 5040 36252 5046 36304
rect 750 36184 756 36236
rect 808 36224 814 36236
rect 1118 36224 1124 36236
rect 808 36196 1124 36224
rect 808 36184 814 36196
rect 1118 36184 1124 36196
rect 1176 36224 1182 36236
rect 1176 36196 2774 36224
rect 1176 36184 1182 36196
rect 1949 36159 2007 36165
rect 1949 36125 1961 36159
rect 1995 36156 2007 36159
rect 2133 36159 2191 36165
rect 1995 36128 2084 36156
rect 1995 36125 2007 36128
rect 1949 36119 2007 36125
rect 2056 36020 2084 36128
rect 2133 36125 2145 36159
rect 2179 36125 2191 36159
rect 2746 36156 2774 36196
rect 3053 36159 3111 36165
rect 3053 36156 3065 36159
rect 2746 36128 3065 36156
rect 2133 36119 2191 36125
rect 3053 36125 3065 36128
rect 3099 36125 3111 36159
rect 3053 36119 3111 36125
rect 3237 36159 3295 36165
rect 3237 36125 3249 36159
rect 3283 36156 3295 36159
rect 3970 36156 3976 36168
rect 3283 36128 3976 36156
rect 3283 36125 3295 36128
rect 3237 36119 3295 36125
rect 2148 36088 2176 36119
rect 3970 36116 3976 36128
rect 4028 36116 4034 36168
rect 9858 36156 9864 36168
rect 9819 36128 9864 36156
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 3602 36088 3608 36100
rect 2148 36060 3608 36088
rect 3602 36048 3608 36060
rect 3660 36048 3666 36100
rect 2958 36020 2964 36032
rect 2056 35992 2964 36020
rect 2958 35980 2964 35992
rect 3016 35980 3022 36032
rect 10042 36020 10048 36032
rect 10003 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 1104 35930 10856 35952
rect 1104 35878 4213 35930
rect 4265 35878 4277 35930
rect 4329 35878 4341 35930
rect 4393 35878 4405 35930
rect 4457 35878 4469 35930
rect 4521 35878 7477 35930
rect 7529 35878 7541 35930
rect 7593 35878 7605 35930
rect 7657 35878 7669 35930
rect 7721 35878 7733 35930
rect 7785 35878 10856 35930
rect 1104 35856 10856 35878
rect 2317 35819 2375 35825
rect 2317 35785 2329 35819
rect 2363 35816 2375 35819
rect 4706 35816 4712 35828
rect 2363 35788 4712 35816
rect 2363 35785 2375 35788
rect 2317 35779 2375 35785
rect 4706 35776 4712 35788
rect 4764 35776 4770 35828
rect 2133 35683 2191 35689
rect 2133 35649 2145 35683
rect 2179 35649 2191 35683
rect 2314 35680 2320 35692
rect 2275 35652 2320 35680
rect 2133 35643 2191 35649
rect 2148 35612 2176 35643
rect 2314 35640 2320 35652
rect 2372 35640 2378 35692
rect 2869 35683 2927 35689
rect 2869 35649 2881 35683
rect 2915 35680 2927 35683
rect 3694 35680 3700 35692
rect 2915 35652 3700 35680
rect 2915 35649 2927 35652
rect 2869 35643 2927 35649
rect 3694 35640 3700 35652
rect 3752 35640 3758 35692
rect 2958 35612 2964 35624
rect 2148 35584 2964 35612
rect 2958 35572 2964 35584
rect 3016 35572 3022 35624
rect 3050 35544 3056 35556
rect 3011 35516 3056 35544
rect 3050 35504 3056 35516
rect 3108 35504 3114 35556
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5845 35386
rect 5897 35334 5909 35386
rect 5961 35334 5973 35386
rect 6025 35334 6037 35386
rect 6089 35334 6101 35386
rect 6153 35334 9109 35386
rect 9161 35334 9173 35386
rect 9225 35334 9237 35386
rect 9289 35334 9301 35386
rect 9353 35334 9365 35386
rect 9417 35334 10856 35386
rect 1104 35312 10856 35334
rect 3973 35275 4031 35281
rect 3973 35241 3985 35275
rect 4019 35272 4031 35275
rect 9858 35272 9864 35284
rect 4019 35244 9864 35272
rect 4019 35241 4031 35244
rect 3973 35235 4031 35241
rect 9858 35232 9864 35244
rect 9916 35232 9922 35284
rect 2777 35207 2835 35213
rect 2777 35173 2789 35207
rect 2823 35204 2835 35207
rect 8846 35204 8852 35216
rect 2823 35176 8852 35204
rect 2823 35173 2835 35176
rect 2777 35167 2835 35173
rect 8846 35164 8852 35176
rect 8904 35164 8910 35216
rect 1949 35071 2007 35077
rect 1949 35037 1961 35071
rect 1995 35068 2007 35071
rect 1995 35040 2084 35068
rect 1995 35037 2007 35040
rect 1949 35031 2007 35037
rect 2056 34932 2084 35040
rect 2130 35028 2136 35080
rect 2188 35068 2194 35080
rect 2777 35071 2835 35077
rect 2777 35068 2789 35071
rect 2188 35040 2789 35068
rect 2188 35028 2194 35040
rect 2777 35037 2789 35040
rect 2823 35068 2835 35071
rect 2958 35068 2964 35080
rect 2823 35040 2964 35068
rect 2823 35037 2835 35040
rect 2777 35031 2835 35037
rect 2958 35028 2964 35040
rect 3016 35028 3022 35080
rect 3053 35071 3111 35077
rect 3053 35037 3065 35071
rect 3099 35068 3111 35071
rect 3602 35068 3608 35080
rect 3099 35040 3608 35068
rect 3099 35037 3111 35040
rect 3053 35031 3111 35037
rect 3602 35028 3608 35040
rect 3660 35068 3666 35080
rect 3789 35071 3847 35077
rect 3789 35068 3801 35071
rect 3660 35040 3801 35068
rect 3660 35028 3666 35040
rect 3789 35037 3801 35040
rect 3835 35037 3847 35071
rect 3970 35068 3976 35080
rect 3931 35040 3976 35068
rect 3789 35031 3847 35037
rect 3970 35028 3976 35040
rect 4028 35028 4034 35080
rect 9858 35068 9864 35080
rect 9819 35040 9864 35068
rect 9858 35028 9864 35040
rect 9916 35028 9922 35080
rect 2225 35003 2283 35009
rect 2225 34969 2237 35003
rect 2271 35000 2283 35003
rect 5442 35000 5448 35012
rect 2271 34972 5448 35000
rect 2271 34969 2283 34972
rect 2225 34963 2283 34969
rect 5442 34960 5448 34972
rect 5500 34960 5506 35012
rect 2958 34932 2964 34944
rect 2056 34904 2964 34932
rect 2958 34892 2964 34904
rect 3016 34892 3022 34944
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 1104 34842 10856 34864
rect 1104 34790 4213 34842
rect 4265 34790 4277 34842
rect 4329 34790 4341 34842
rect 4393 34790 4405 34842
rect 4457 34790 4469 34842
rect 4521 34790 7477 34842
rect 7529 34790 7541 34842
rect 7593 34790 7605 34842
rect 7657 34790 7669 34842
rect 7721 34790 7733 34842
rect 7785 34790 10856 34842
rect 1104 34768 10856 34790
rect 3050 34728 3056 34740
rect 1688 34700 3056 34728
rect 1688 34660 1716 34700
rect 3050 34688 3056 34700
rect 3108 34688 3114 34740
rect 3234 34728 3240 34740
rect 3195 34700 3240 34728
rect 3234 34688 3240 34700
rect 3292 34688 3298 34740
rect 1596 34632 1716 34660
rect 1857 34663 1915 34669
rect 1596 34601 1624 34632
rect 1857 34629 1869 34663
rect 1903 34660 1915 34663
rect 8754 34660 8760 34672
rect 1903 34632 8760 34660
rect 1903 34629 1915 34632
rect 1857 34623 1915 34629
rect 8754 34620 8760 34632
rect 8812 34620 8818 34672
rect 1581 34595 1639 34601
rect 1581 34561 1593 34595
rect 1627 34561 1639 34595
rect 1581 34555 1639 34561
rect 1673 34595 1731 34601
rect 1673 34561 1685 34595
rect 1719 34592 1731 34595
rect 2130 34592 2136 34604
rect 1719 34564 2136 34592
rect 1719 34561 1731 34564
rect 1673 34555 1731 34561
rect 845 34527 903 34533
rect 845 34493 857 34527
rect 891 34524 903 34527
rect 1688 34524 1716 34555
rect 2130 34552 2136 34564
rect 2188 34552 2194 34604
rect 2406 34552 2412 34604
rect 2464 34592 2470 34604
rect 2593 34595 2651 34601
rect 2593 34592 2605 34595
rect 2464 34564 2605 34592
rect 2464 34552 2470 34564
rect 2593 34561 2605 34564
rect 2639 34561 2651 34595
rect 2593 34555 2651 34561
rect 3053 34595 3111 34601
rect 3053 34561 3065 34595
rect 3099 34592 3111 34595
rect 3142 34592 3148 34604
rect 3099 34564 3148 34592
rect 3099 34561 3111 34564
rect 3053 34555 3111 34561
rect 3142 34552 3148 34564
rect 3200 34552 3206 34604
rect 9674 34552 9680 34604
rect 9732 34592 9738 34604
rect 9861 34595 9919 34601
rect 9861 34592 9873 34595
rect 9732 34564 9873 34592
rect 9732 34552 9738 34564
rect 9861 34561 9873 34564
rect 9907 34561 9919 34595
rect 9861 34555 9919 34561
rect 891 34496 1716 34524
rect 891 34493 903 34496
rect 845 34487 903 34493
rect 2130 34416 2136 34468
rect 2188 34456 2194 34468
rect 11241 34459 11299 34465
rect 11241 34456 11253 34459
rect 2188 34428 11253 34456
rect 2188 34416 2194 34428
rect 11241 34425 11253 34428
rect 11287 34425 11299 34459
rect 11241 34419 11299 34425
rect 2406 34388 2412 34400
rect 2367 34360 2412 34388
rect 2406 34348 2412 34360
rect 2464 34348 2470 34400
rect 10042 34388 10048 34400
rect 10003 34360 10048 34388
rect 10042 34348 10048 34360
rect 10100 34348 10106 34400
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5845 34298
rect 5897 34246 5909 34298
rect 5961 34246 5973 34298
rect 6025 34246 6037 34298
rect 6089 34246 6101 34298
rect 6153 34246 9109 34298
rect 9161 34246 9173 34298
rect 9225 34246 9237 34298
rect 9289 34246 9301 34298
rect 9353 34246 9365 34298
rect 9417 34246 10856 34298
rect 1104 34224 10856 34246
rect 1486 34184 1492 34196
rect 1447 34156 1492 34184
rect 1486 34144 1492 34156
rect 1544 34144 1550 34196
rect 3053 34187 3111 34193
rect 1688 34156 3004 34184
rect 1688 33989 1716 34156
rect 2976 34116 3004 34156
rect 3053 34153 3065 34187
rect 3099 34184 3111 34187
rect 9766 34184 9772 34196
rect 3099 34156 9772 34184
rect 3099 34153 3111 34156
rect 3053 34147 3111 34153
rect 9766 34144 9772 34156
rect 9824 34144 9830 34196
rect 8570 34116 8576 34128
rect 2976 34088 8576 34116
rect 8570 34076 8576 34088
rect 8628 34076 8634 34128
rect 1673 33983 1731 33989
rect 1673 33949 1685 33983
rect 1719 33949 1731 33983
rect 2130 33980 2136 33992
rect 2091 33952 2136 33980
rect 1673 33943 1731 33949
rect 2130 33940 2136 33952
rect 2188 33940 2194 33992
rect 2869 33983 2927 33989
rect 2869 33949 2881 33983
rect 2915 33949 2927 33983
rect 2869 33943 2927 33949
rect 3053 33983 3111 33989
rect 3053 33949 3065 33983
rect 3099 33980 3111 33983
rect 3234 33980 3240 33992
rect 3099 33952 3240 33980
rect 3099 33949 3111 33952
rect 3053 33943 3111 33949
rect 2884 33912 2912 33943
rect 3234 33940 3240 33952
rect 3292 33980 3298 33992
rect 3970 33980 3976 33992
rect 3292 33952 3976 33980
rect 3292 33940 3298 33952
rect 3970 33940 3976 33952
rect 4028 33940 4034 33992
rect 4614 33912 4620 33924
rect 2884 33884 4620 33912
rect 3068 33856 3096 33884
rect 4614 33872 4620 33884
rect 4672 33872 4678 33924
rect 2314 33844 2320 33856
rect 2275 33816 2320 33844
rect 2314 33804 2320 33816
rect 2372 33804 2378 33856
rect 3050 33804 3056 33856
rect 3108 33804 3114 33856
rect 1104 33754 10856 33776
rect 1104 33702 4213 33754
rect 4265 33702 4277 33754
rect 4329 33702 4341 33754
rect 4393 33702 4405 33754
rect 4457 33702 4469 33754
rect 4521 33702 7477 33754
rect 7529 33702 7541 33754
rect 7593 33702 7605 33754
rect 7657 33702 7669 33754
rect 7721 33702 7733 33754
rect 7785 33702 10856 33754
rect 1104 33680 10856 33702
rect 2961 33643 3019 33649
rect 2961 33609 2973 33643
rect 3007 33640 3019 33643
rect 3510 33640 3516 33652
rect 3007 33612 3516 33640
rect 3007 33609 3019 33612
rect 2961 33603 3019 33609
rect 3510 33600 3516 33612
rect 3568 33600 3574 33652
rect 1397 33507 1455 33513
rect 1397 33473 1409 33507
rect 1443 33504 1455 33507
rect 1578 33504 1584 33516
rect 1443 33476 1584 33504
rect 1443 33473 1455 33476
rect 1397 33467 1455 33473
rect 1578 33464 1584 33476
rect 1636 33464 1642 33516
rect 2038 33464 2044 33516
rect 2096 33504 2102 33516
rect 2133 33507 2191 33513
rect 2133 33504 2145 33507
rect 2096 33476 2145 33504
rect 2096 33464 2102 33476
rect 2133 33473 2145 33476
rect 2179 33473 2191 33507
rect 2133 33467 2191 33473
rect 2869 33507 2927 33513
rect 2869 33473 2881 33507
rect 2915 33504 2927 33507
rect 3418 33504 3424 33516
rect 2915 33476 3424 33504
rect 2915 33473 2927 33476
rect 2869 33467 2927 33473
rect 3418 33464 3424 33476
rect 3476 33464 3482 33516
rect 9766 33464 9772 33516
rect 9824 33504 9830 33516
rect 9861 33507 9919 33513
rect 9861 33504 9873 33507
rect 9824 33476 9873 33504
rect 9824 33464 9830 33476
rect 9861 33473 9873 33476
rect 9907 33473 9919 33507
rect 9861 33467 9919 33473
rect 2130 33328 2136 33380
rect 2188 33368 2194 33380
rect 3326 33368 3332 33380
rect 2188 33340 3332 33368
rect 2188 33328 2194 33340
rect 3326 33328 3332 33340
rect 3384 33328 3390 33380
rect 10042 33368 10048 33380
rect 10003 33340 10048 33368
rect 10042 33328 10048 33340
rect 10100 33328 10106 33380
rect 1486 33260 1492 33312
rect 1544 33300 1550 33312
rect 1581 33303 1639 33309
rect 1581 33300 1593 33303
rect 1544 33272 1593 33300
rect 1544 33260 1550 33272
rect 1581 33269 1593 33272
rect 1627 33269 1639 33303
rect 2314 33300 2320 33312
rect 2275 33272 2320 33300
rect 1581 33263 1639 33269
rect 2314 33260 2320 33272
rect 2372 33260 2378 33312
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5845 33210
rect 5897 33158 5909 33210
rect 5961 33158 5973 33210
rect 6025 33158 6037 33210
rect 6089 33158 6101 33210
rect 6153 33158 9109 33210
rect 9161 33158 9173 33210
rect 9225 33158 9237 33210
rect 9289 33158 9301 33210
rect 9353 33158 9365 33210
rect 9417 33158 10856 33210
rect 1104 33136 10856 33158
rect 3973 33099 4031 33105
rect 3973 33065 3985 33099
rect 4019 33096 4031 33099
rect 9858 33096 9864 33108
rect 4019 33068 9864 33096
rect 4019 33065 4031 33068
rect 3973 33059 4031 33065
rect 9858 33056 9864 33068
rect 9916 33056 9922 33108
rect 3053 33031 3111 33037
rect 3053 32997 3065 33031
rect 3099 33028 3111 33031
rect 9674 33028 9680 33040
rect 3099 33000 9680 33028
rect 3099 32997 3111 33000
rect 3053 32991 3111 32997
rect 9674 32988 9680 33000
rect 9732 32988 9738 33040
rect 3252 32932 4016 32960
rect 3252 32904 3280 32932
rect 1394 32892 1400 32904
rect 1355 32864 1400 32892
rect 1394 32852 1400 32864
rect 1452 32852 1458 32904
rect 1946 32852 1952 32904
rect 2004 32892 2010 32904
rect 2133 32895 2191 32901
rect 2133 32892 2145 32895
rect 2004 32864 2145 32892
rect 2004 32852 2010 32864
rect 2133 32861 2145 32864
rect 2179 32861 2191 32895
rect 2133 32855 2191 32861
rect 2869 32895 2927 32901
rect 2869 32861 2881 32895
rect 2915 32892 2927 32895
rect 2958 32892 2964 32904
rect 2915 32864 2964 32892
rect 2915 32861 2927 32864
rect 2869 32855 2927 32861
rect 2958 32852 2964 32864
rect 3016 32852 3022 32904
rect 3053 32895 3111 32901
rect 3053 32861 3065 32895
rect 3099 32892 3111 32895
rect 3234 32892 3240 32904
rect 3099 32864 3240 32892
rect 3099 32861 3111 32864
rect 3053 32855 3111 32861
rect 3234 32852 3240 32864
rect 3292 32852 3298 32904
rect 3694 32852 3700 32904
rect 3752 32892 3758 32904
rect 3988 32901 4016 32932
rect 3789 32895 3847 32901
rect 3789 32892 3801 32895
rect 3752 32864 3801 32892
rect 3752 32852 3758 32864
rect 3789 32861 3801 32864
rect 3835 32861 3847 32895
rect 3789 32855 3847 32861
rect 3973 32895 4031 32901
rect 3973 32861 3985 32895
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 9861 32895 9919 32901
rect 9861 32861 9873 32895
rect 9907 32892 9919 32895
rect 11149 32895 11207 32901
rect 11149 32892 11161 32895
rect 9907 32864 11161 32892
rect 9907 32861 9919 32864
rect 9861 32855 9919 32861
rect 11149 32861 11161 32864
rect 11195 32861 11207 32895
rect 11149 32855 11207 32861
rect 3804 32824 3832 32855
rect 4062 32824 4068 32836
rect 3804 32796 4068 32824
rect 4062 32784 4068 32796
rect 4120 32784 4126 32836
rect 1578 32756 1584 32768
rect 1539 32728 1584 32756
rect 1578 32716 1584 32728
rect 1636 32716 1642 32768
rect 1670 32716 1676 32768
rect 1728 32756 1734 32768
rect 1946 32756 1952 32768
rect 1728 32728 1952 32756
rect 1728 32716 1734 32728
rect 1946 32716 1952 32728
rect 2004 32716 2010 32768
rect 2314 32756 2320 32768
rect 2275 32728 2320 32756
rect 2314 32716 2320 32728
rect 2372 32716 2378 32768
rect 3694 32716 3700 32768
rect 3752 32756 3758 32768
rect 3878 32756 3884 32768
rect 3752 32728 3884 32756
rect 3752 32716 3758 32728
rect 3878 32716 3884 32728
rect 3936 32716 3942 32768
rect 10042 32756 10048 32768
rect 10003 32728 10048 32756
rect 10042 32716 10048 32728
rect 10100 32716 10106 32768
rect 1104 32666 10856 32688
rect 1104 32614 4213 32666
rect 4265 32614 4277 32666
rect 4329 32614 4341 32666
rect 4393 32614 4405 32666
rect 4457 32614 4469 32666
rect 4521 32614 7477 32666
rect 7529 32614 7541 32666
rect 7593 32614 7605 32666
rect 7657 32614 7669 32666
rect 7721 32614 7733 32666
rect 7785 32614 10856 32666
rect 1104 32592 10856 32614
rect 2869 32555 2927 32561
rect 2869 32521 2881 32555
rect 2915 32552 2927 32555
rect 9766 32552 9772 32564
rect 2915 32524 9772 32552
rect 2915 32521 2927 32524
rect 2869 32515 2927 32521
rect 9766 32512 9772 32524
rect 9824 32512 9830 32564
rect 3970 32484 3976 32496
rect 1688 32456 3976 32484
rect 1688 32425 1716 32456
rect 3970 32444 3976 32456
rect 4028 32444 4034 32496
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32385 1731 32419
rect 1673 32379 1731 32385
rect 2038 32376 2044 32428
rect 2096 32416 2102 32428
rect 2406 32416 2412 32428
rect 2096 32388 2412 32416
rect 2096 32376 2102 32388
rect 2406 32376 2412 32388
rect 2464 32416 2470 32428
rect 2777 32419 2835 32425
rect 2777 32416 2789 32419
rect 2464 32388 2789 32416
rect 2464 32376 2470 32388
rect 2777 32385 2789 32388
rect 2823 32385 2835 32419
rect 2777 32379 2835 32385
rect 2961 32419 3019 32425
rect 2961 32385 2973 32419
rect 3007 32416 3019 32419
rect 3234 32416 3240 32428
rect 3007 32388 3240 32416
rect 3007 32385 3019 32388
rect 2961 32379 3019 32385
rect 3234 32376 3240 32388
rect 3292 32376 3298 32428
rect 937 32351 995 32357
rect 937 32317 949 32351
rect 983 32348 995 32351
rect 1762 32348 1768 32360
rect 983 32320 1768 32348
rect 983 32317 995 32320
rect 937 32311 995 32317
rect 1762 32308 1768 32320
rect 1820 32308 1826 32360
rect 1486 32212 1492 32224
rect 1447 32184 1492 32212
rect 1486 32172 1492 32184
rect 1544 32172 1550 32224
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5845 32122
rect 5897 32070 5909 32122
rect 5961 32070 5973 32122
rect 6025 32070 6037 32122
rect 6089 32070 6101 32122
rect 6153 32070 9109 32122
rect 9161 32070 9173 32122
rect 9225 32070 9237 32122
rect 9289 32070 9301 32122
rect 9353 32070 9365 32122
rect 9417 32070 10856 32122
rect 1104 32048 10856 32070
rect 2041 32011 2099 32017
rect 2041 31977 2053 32011
rect 2087 32008 2099 32011
rect 5258 32008 5264 32020
rect 2087 31980 5264 32008
rect 2087 31977 2099 31980
rect 2041 31971 2099 31977
rect 5258 31968 5264 31980
rect 5316 31968 5322 32020
rect 2685 31943 2743 31949
rect 2685 31909 2697 31943
rect 2731 31940 2743 31943
rect 2774 31940 2780 31952
rect 2731 31912 2780 31940
rect 2731 31909 2743 31912
rect 2685 31903 2743 31909
rect 2774 31900 2780 31912
rect 2832 31900 2838 31952
rect 10042 31940 10048 31952
rect 10003 31912 10048 31940
rect 10042 31900 10048 31912
rect 10100 31900 10106 31952
rect 3786 31872 3792 31884
rect 2056 31844 3792 31872
rect 2056 31813 2084 31844
rect 3786 31832 3792 31844
rect 3844 31832 3850 31884
rect 2041 31807 2099 31813
rect 2041 31773 2053 31807
rect 2087 31773 2099 31807
rect 2498 31804 2504 31816
rect 2459 31776 2504 31804
rect 2041 31767 2099 31773
rect 2498 31764 2504 31776
rect 2556 31764 2562 31816
rect 9861 31807 9919 31813
rect 9861 31773 9873 31807
rect 9907 31804 9919 31807
rect 11241 31807 11299 31813
rect 11241 31804 11253 31807
rect 9907 31776 11253 31804
rect 9907 31773 9919 31776
rect 9861 31767 9919 31773
rect 11241 31773 11253 31776
rect 11287 31773 11299 31807
rect 11241 31767 11299 31773
rect 2498 31628 2504 31680
rect 2556 31668 2562 31680
rect 3142 31668 3148 31680
rect 2556 31640 3148 31668
rect 2556 31628 2562 31640
rect 3142 31628 3148 31640
rect 3200 31628 3206 31680
rect 1104 31578 10856 31600
rect 1104 31526 4213 31578
rect 4265 31526 4277 31578
rect 4329 31526 4341 31578
rect 4393 31526 4405 31578
rect 4457 31526 4469 31578
rect 4521 31526 7477 31578
rect 7529 31526 7541 31578
rect 7593 31526 7605 31578
rect 7657 31526 7669 31578
rect 7721 31526 7733 31578
rect 7785 31526 10856 31578
rect 1104 31504 10856 31526
rect 2409 31467 2467 31473
rect 2409 31433 2421 31467
rect 2455 31464 2467 31467
rect 6638 31464 6644 31476
rect 2455 31436 6644 31464
rect 2455 31433 2467 31436
rect 2409 31427 2467 31433
rect 6638 31424 6644 31436
rect 6696 31424 6702 31476
rect 290 31356 296 31408
rect 348 31396 354 31408
rect 1581 31399 1639 31405
rect 1581 31396 1593 31399
rect 348 31368 1593 31396
rect 348 31356 354 31368
rect 1581 31365 1593 31368
rect 1627 31365 1639 31399
rect 1581 31359 1639 31365
rect 1857 31331 1915 31337
rect 1857 31297 1869 31331
rect 1903 31297 1915 31331
rect 1857 31291 1915 31297
rect 2593 31331 2651 31337
rect 2593 31297 2605 31331
rect 2639 31328 2651 31331
rect 3050 31328 3056 31340
rect 2639 31300 3056 31328
rect 2639 31297 2651 31300
rect 2593 31291 2651 31297
rect 1872 31260 1900 31291
rect 3050 31288 3056 31300
rect 3108 31288 3114 31340
rect 9861 31331 9919 31337
rect 9861 31297 9873 31331
rect 9907 31328 9919 31331
rect 11057 31331 11115 31337
rect 11057 31328 11069 31331
rect 9907 31300 11069 31328
rect 9907 31297 9919 31300
rect 9861 31291 9919 31297
rect 11057 31297 11069 31300
rect 11103 31297 11115 31331
rect 11057 31291 11115 31297
rect 3418 31260 3424 31272
rect 1872 31232 3424 31260
rect 3418 31220 3424 31232
rect 3476 31220 3482 31272
rect 2130 31084 2136 31136
rect 2188 31124 2194 31136
rect 2406 31124 2412 31136
rect 2188 31096 2412 31124
rect 2188 31084 2194 31096
rect 2406 31084 2412 31096
rect 2464 31084 2470 31136
rect 10042 31124 10048 31136
rect 10003 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5845 31034
rect 5897 30982 5909 31034
rect 5961 30982 5973 31034
rect 6025 30982 6037 31034
rect 6089 30982 6101 31034
rect 6153 30982 9109 31034
rect 9161 30982 9173 31034
rect 9225 30982 9237 31034
rect 9289 30982 9301 31034
rect 9353 30982 9365 31034
rect 9417 30982 10856 31034
rect 1104 30960 10856 30982
rect 382 30880 388 30932
rect 440 30920 446 30932
rect 2041 30923 2099 30929
rect 2041 30920 2053 30923
rect 440 30892 2053 30920
rect 440 30880 446 30892
rect 2041 30889 2053 30892
rect 2087 30889 2099 30923
rect 2041 30883 2099 30889
rect 2777 30923 2835 30929
rect 2777 30889 2789 30923
rect 2823 30920 2835 30923
rect 3510 30920 3516 30932
rect 2823 30892 3516 30920
rect 2823 30889 2835 30892
rect 2777 30883 2835 30889
rect 3510 30880 3516 30892
rect 3568 30880 3574 30932
rect 3786 30920 3792 30932
rect 3747 30892 3792 30920
rect 3786 30880 3792 30892
rect 3844 30880 3850 30932
rect 1670 30812 1676 30864
rect 1728 30852 1734 30864
rect 8662 30852 8668 30864
rect 1728 30824 8668 30852
rect 1728 30812 1734 30824
rect 8662 30812 8668 30824
rect 8720 30812 8726 30864
rect 2590 30744 2596 30796
rect 2648 30784 2654 30796
rect 7098 30784 7104 30796
rect 2648 30756 7104 30784
rect 2648 30744 2654 30756
rect 7098 30744 7104 30756
rect 7156 30744 7162 30796
rect 2225 30719 2283 30725
rect 2225 30685 2237 30719
rect 2271 30685 2283 30719
rect 2225 30679 2283 30685
rect 2869 30719 2927 30725
rect 2869 30685 2881 30719
rect 2915 30716 2927 30719
rect 3510 30716 3516 30728
rect 2915 30688 3516 30716
rect 2915 30685 2927 30688
rect 2869 30679 2927 30685
rect 2240 30648 2268 30679
rect 3510 30676 3516 30688
rect 3568 30676 3574 30728
rect 3970 30716 3976 30728
rect 3931 30688 3976 30716
rect 3970 30676 3976 30688
rect 4028 30676 4034 30728
rect 9401 30719 9459 30725
rect 9401 30685 9413 30719
rect 9447 30716 9459 30719
rect 9490 30716 9496 30728
rect 9447 30688 9496 30716
rect 9447 30685 9459 30688
rect 9401 30679 9459 30685
rect 9490 30676 9496 30688
rect 9548 30676 9554 30728
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30716 9919 30719
rect 10965 30719 11023 30725
rect 10965 30716 10977 30719
rect 9907 30688 10977 30716
rect 9907 30685 9919 30688
rect 9861 30679 9919 30685
rect 10965 30685 10977 30688
rect 11011 30685 11023 30719
rect 10965 30679 11023 30685
rect 2958 30648 2964 30660
rect 2240 30620 2964 30648
rect 2958 30608 2964 30620
rect 3016 30608 3022 30660
rect 10042 30580 10048 30592
rect 10003 30552 10048 30580
rect 10042 30540 10048 30552
rect 10100 30540 10106 30592
rect 1104 30490 10856 30512
rect 1104 30438 4213 30490
rect 4265 30438 4277 30490
rect 4329 30438 4341 30490
rect 4393 30438 4405 30490
rect 4457 30438 4469 30490
rect 4521 30438 7477 30490
rect 7529 30438 7541 30490
rect 7593 30438 7605 30490
rect 7657 30438 7669 30490
rect 7721 30438 7733 30490
rect 7785 30438 10856 30490
rect 1104 30416 10856 30438
rect 2409 30379 2467 30385
rect 2409 30345 2421 30379
rect 2455 30345 2467 30379
rect 2409 30339 2467 30345
rect 845 30311 903 30317
rect 845 30277 857 30311
rect 891 30308 903 30311
rect 2424 30308 2452 30339
rect 3142 30336 3148 30388
rect 3200 30376 3206 30388
rect 3697 30379 3755 30385
rect 3697 30376 3709 30379
rect 3200 30348 3709 30376
rect 3200 30336 3206 30348
rect 3697 30345 3709 30348
rect 3743 30345 3755 30379
rect 3697 30339 3755 30345
rect 2590 30308 2596 30320
rect 891 30280 2268 30308
rect 2424 30280 2596 30308
rect 891 30277 903 30280
rect 845 30271 903 30277
rect 2240 30252 2268 30280
rect 2590 30268 2596 30280
rect 2648 30268 2654 30320
rect 5350 30308 5356 30320
rect 3804 30280 5356 30308
rect 1670 30240 1676 30252
rect 1631 30212 1676 30240
rect 1670 30200 1676 30212
rect 1728 30200 1734 30252
rect 2222 30240 2228 30252
rect 2183 30212 2228 30240
rect 2222 30200 2228 30212
rect 2280 30200 2286 30252
rect 2409 30243 2467 30249
rect 2409 30209 2421 30243
rect 2455 30209 2467 30243
rect 2409 30203 2467 30209
rect 3053 30243 3111 30249
rect 3053 30209 3065 30243
rect 3099 30209 3111 30243
rect 3053 30203 3111 30209
rect 3237 30243 3295 30249
rect 3237 30209 3249 30243
rect 3283 30240 3295 30243
rect 3804 30240 3832 30280
rect 5350 30268 5356 30280
rect 5408 30268 5414 30320
rect 3283 30212 3832 30240
rect 3881 30243 3939 30249
rect 3283 30209 3295 30212
rect 3237 30203 3295 30209
rect 3881 30209 3893 30243
rect 3927 30209 3939 30243
rect 3881 30203 3939 30209
rect 2130 30132 2136 30184
rect 2188 30172 2194 30184
rect 2424 30172 2452 30203
rect 2188 30144 2452 30172
rect 2188 30132 2194 30144
rect 1486 30104 1492 30116
rect 1447 30076 1492 30104
rect 1486 30064 1492 30076
rect 1544 30064 1550 30116
rect 3068 30048 3096 30203
rect 3896 30116 3924 30203
rect 3878 30064 3884 30116
rect 3936 30064 3942 30116
rect 3050 29996 3056 30048
rect 3108 29996 3114 30048
rect 10134 30036 10140 30048
rect 10095 30008 10140 30036
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5845 29946
rect 5897 29894 5909 29946
rect 5961 29894 5973 29946
rect 6025 29894 6037 29946
rect 6089 29894 6101 29946
rect 6153 29894 9109 29946
rect 9161 29894 9173 29946
rect 9225 29894 9237 29946
rect 9289 29894 9301 29946
rect 9353 29894 9365 29946
rect 9417 29894 10856 29946
rect 1104 29872 10856 29894
rect 106 29792 112 29844
rect 164 29832 170 29844
rect 1489 29835 1547 29841
rect 1489 29832 1501 29835
rect 164 29804 1501 29832
rect 164 29792 170 29804
rect 1489 29801 1501 29804
rect 1535 29801 1547 29835
rect 1489 29795 1547 29801
rect 3418 29792 3424 29844
rect 3476 29832 3482 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 3476 29804 3801 29832
rect 3476 29792 3482 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 3789 29795 3847 29801
rect 2130 29724 2136 29776
rect 2188 29764 2194 29776
rect 3237 29767 3295 29773
rect 2188 29736 2774 29764
rect 2188 29724 2194 29736
rect 1302 29656 1308 29708
rect 1360 29696 1366 29708
rect 2225 29699 2283 29705
rect 2225 29696 2237 29699
rect 1360 29668 2237 29696
rect 1360 29656 1366 29668
rect 2225 29665 2237 29668
rect 2271 29665 2283 29699
rect 2225 29659 2283 29665
rect 1578 29628 1584 29640
rect 1539 29600 1584 29628
rect 1578 29588 1584 29600
rect 1636 29588 1642 29640
rect 2317 29631 2375 29637
rect 2317 29597 2329 29631
rect 2363 29597 2375 29631
rect 2317 29591 2375 29597
rect 2593 29631 2651 29637
rect 2593 29597 2605 29631
rect 2639 29597 2651 29631
rect 2746 29628 2774 29736
rect 3237 29733 3249 29767
rect 3283 29764 3295 29767
rect 11149 29767 11207 29773
rect 11149 29764 11161 29767
rect 3283 29736 11161 29764
rect 3283 29733 3295 29736
rect 3237 29727 3295 29733
rect 11149 29733 11161 29736
rect 11195 29733 11207 29767
rect 11149 29727 11207 29733
rect 3053 29631 3111 29637
rect 3053 29628 3065 29631
rect 2746 29600 3065 29628
rect 2593 29591 2651 29597
rect 3053 29597 3065 29600
rect 3099 29597 3111 29631
rect 3053 29591 3111 29597
rect 474 29520 480 29572
rect 532 29560 538 29572
rect 1762 29560 1768 29572
rect 532 29532 1768 29560
rect 532 29520 538 29532
rect 1762 29520 1768 29532
rect 1820 29560 1826 29572
rect 2332 29560 2360 29591
rect 1820 29532 2360 29560
rect 2608 29560 2636 29591
rect 3234 29588 3240 29640
rect 3292 29628 3298 29640
rect 3418 29628 3424 29640
rect 3292 29600 3424 29628
rect 3292 29588 3298 29600
rect 3418 29588 3424 29600
rect 3476 29588 3482 29640
rect 3970 29628 3976 29640
rect 3931 29600 3976 29628
rect 3970 29588 3976 29600
rect 4028 29588 4034 29640
rect 4706 29560 4712 29572
rect 2608 29532 4712 29560
rect 1820 29520 1826 29532
rect 4706 29520 4712 29532
rect 4764 29520 4770 29572
rect 3878 29452 3884 29504
rect 3936 29492 3942 29504
rect 4614 29492 4620 29504
rect 3936 29464 4620 29492
rect 3936 29452 3942 29464
rect 4614 29452 4620 29464
rect 4672 29452 4678 29504
rect 1104 29402 10856 29424
rect 1104 29350 4213 29402
rect 4265 29350 4277 29402
rect 4329 29350 4341 29402
rect 4393 29350 4405 29402
rect 4457 29350 4469 29402
rect 4521 29350 7477 29402
rect 7529 29350 7541 29402
rect 7593 29350 7605 29402
rect 7657 29350 7669 29402
rect 7721 29350 7733 29402
rect 7785 29350 10856 29402
rect 1104 29328 10856 29350
rect 1578 29288 1584 29300
rect 1539 29260 1584 29288
rect 1578 29248 1584 29260
rect 1636 29248 1642 29300
rect 2501 29291 2559 29297
rect 2501 29257 2513 29291
rect 2547 29288 2559 29291
rect 2547 29260 2774 29288
rect 2547 29257 2559 29260
rect 2501 29251 2559 29257
rect 1302 29180 1308 29232
rect 1360 29220 1366 29232
rect 2746 29220 2774 29260
rect 2958 29248 2964 29300
rect 3016 29288 3022 29300
rect 3053 29291 3111 29297
rect 3053 29288 3065 29291
rect 3016 29260 3065 29288
rect 3016 29248 3022 29260
rect 3053 29257 3065 29260
rect 3099 29257 3111 29291
rect 3053 29251 3111 29257
rect 5074 29220 5080 29232
rect 1360 29192 2544 29220
rect 2746 29192 5080 29220
rect 1360 29180 1366 29192
rect 1394 29152 1400 29164
rect 1355 29124 1400 29152
rect 1394 29112 1400 29124
rect 1452 29112 1458 29164
rect 1578 29112 1584 29164
rect 1636 29152 1642 29164
rect 2130 29152 2136 29164
rect 1636 29124 2136 29152
rect 1636 29112 1642 29124
rect 2130 29112 2136 29124
rect 2188 29112 2194 29164
rect 2516 29161 2544 29192
rect 5074 29180 5080 29192
rect 5132 29180 5138 29232
rect 2317 29155 2375 29161
rect 2317 29121 2329 29155
rect 2363 29121 2375 29155
rect 2317 29115 2375 29121
rect 2501 29155 2559 29161
rect 2501 29121 2513 29155
rect 2547 29121 2559 29155
rect 3234 29152 3240 29164
rect 3195 29124 3240 29152
rect 2501 29115 2559 29121
rect 1762 29044 1768 29096
rect 1820 29084 1826 29096
rect 2332 29084 2360 29115
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 1820 29056 2360 29084
rect 1820 29044 1826 29056
rect 2148 29028 2176 29056
rect 753 29019 811 29025
rect 753 28985 765 29019
rect 799 29016 811 29019
rect 799 28988 1348 29016
rect 799 28985 811 28988
rect 753 28979 811 28985
rect 937 28951 995 28957
rect 937 28917 949 28951
rect 983 28948 995 28951
rect 1320 28948 1348 28988
rect 2130 28976 2136 29028
rect 2188 28976 2194 29028
rect 983 28920 1348 28948
rect 983 28917 995 28920
rect 937 28911 995 28917
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5845 28858
rect 5897 28806 5909 28858
rect 5961 28806 5973 28858
rect 6025 28806 6037 28858
rect 6089 28806 6101 28858
rect 6153 28806 9109 28858
rect 9161 28806 9173 28858
rect 9225 28806 9237 28858
rect 9289 28806 9301 28858
rect 9353 28806 9365 28858
rect 9417 28806 10856 28858
rect 1104 28784 10856 28806
rect 2314 28744 2320 28756
rect 2275 28716 2320 28744
rect 2314 28704 2320 28716
rect 2372 28704 2378 28756
rect 3050 28744 3056 28756
rect 3011 28716 3056 28744
rect 3050 28704 3056 28716
rect 3108 28704 3114 28756
rect 1765 28679 1823 28685
rect 1765 28645 1777 28679
rect 1811 28676 1823 28679
rect 2498 28676 2504 28688
rect 1811 28648 2504 28676
rect 1811 28645 1823 28648
rect 1765 28639 1823 28645
rect 2498 28636 2504 28648
rect 2556 28636 2562 28688
rect 1762 28540 1768 28552
rect 1723 28512 1768 28540
rect 1762 28500 1768 28512
rect 1820 28500 1826 28552
rect 2409 28543 2467 28549
rect 2409 28509 2421 28543
rect 2455 28509 2467 28543
rect 2866 28540 2872 28552
rect 2827 28512 2872 28540
rect 2409 28503 2467 28509
rect 2424 28472 2452 28503
rect 2866 28500 2872 28512
rect 2924 28500 2930 28552
rect 3234 28472 3240 28484
rect 2424 28444 3240 28472
rect 3234 28432 3240 28444
rect 3292 28432 3298 28484
rect 10134 28404 10140 28416
rect 10095 28376 10140 28404
rect 10134 28364 10140 28376
rect 10192 28364 10198 28416
rect 1104 28314 10856 28336
rect 1104 28262 4213 28314
rect 4265 28262 4277 28314
rect 4329 28262 4341 28314
rect 4393 28262 4405 28314
rect 4457 28262 4469 28314
rect 4521 28262 7477 28314
rect 7529 28262 7541 28314
rect 7593 28262 7605 28314
rect 7657 28262 7669 28314
rect 7721 28262 7733 28314
rect 7785 28262 10856 28314
rect 1104 28240 10856 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 1670 28200 1676 28212
rect 1627 28172 1676 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 1670 28160 1676 28172
rect 1728 28160 1734 28212
rect 1762 28160 1768 28212
rect 1820 28200 1826 28212
rect 2225 28203 2283 28209
rect 2225 28200 2237 28203
rect 1820 28172 2237 28200
rect 1820 28160 1826 28172
rect 2225 28169 2237 28172
rect 2271 28169 2283 28203
rect 2225 28163 2283 28169
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28033 1823 28067
rect 2406 28064 2412 28076
rect 2367 28036 2412 28064
rect 1765 28027 1823 28033
rect 1780 27996 1808 28027
rect 2406 28024 2412 28036
rect 2464 28024 2470 28076
rect 2958 27996 2964 28008
rect 1780 27968 2964 27996
rect 2958 27956 2964 27968
rect 3016 27956 3022 28008
rect 1670 27888 1676 27940
rect 1728 27928 1734 27940
rect 2038 27928 2044 27940
rect 1728 27900 2044 27928
rect 1728 27888 1734 27900
rect 2038 27888 2044 27900
rect 2096 27888 2102 27940
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5845 27770
rect 5897 27718 5909 27770
rect 5961 27718 5973 27770
rect 6025 27718 6037 27770
rect 6089 27718 6101 27770
rect 6153 27718 9109 27770
rect 9161 27718 9173 27770
rect 9225 27718 9237 27770
rect 9289 27718 9301 27770
rect 9353 27718 9365 27770
rect 9417 27718 10856 27770
rect 1104 27696 10856 27718
rect 934 27548 940 27600
rect 992 27588 998 27600
rect 2041 27591 2099 27597
rect 2041 27588 2053 27591
rect 992 27560 2053 27588
rect 992 27548 998 27560
rect 2041 27557 2053 27560
rect 2087 27557 2099 27591
rect 2041 27551 2099 27557
rect 2777 27591 2835 27597
rect 2777 27557 2789 27591
rect 2823 27588 2835 27591
rect 2958 27588 2964 27600
rect 2823 27560 2964 27588
rect 2823 27557 2835 27560
rect 2777 27551 2835 27557
rect 2958 27548 2964 27560
rect 3016 27548 3022 27600
rect 3418 27480 3424 27532
rect 3476 27520 3482 27532
rect 3970 27520 3976 27532
rect 3476 27492 3976 27520
rect 3476 27480 3482 27492
rect 3970 27480 3976 27492
rect 4028 27520 4034 27532
rect 4893 27523 4951 27529
rect 4893 27520 4905 27523
rect 4028 27492 4905 27520
rect 4028 27480 4034 27492
rect 4893 27489 4905 27492
rect 4939 27489 4951 27523
rect 4893 27483 4951 27489
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 2041 27455 2099 27461
rect 2041 27452 2053 27455
rect 1596 27424 2053 27452
rect 1596 27325 1624 27424
rect 2041 27421 2053 27424
rect 2087 27421 2099 27455
rect 2958 27452 2964 27464
rect 2919 27424 2964 27452
rect 2041 27415 2099 27421
rect 2958 27412 2964 27424
rect 3016 27412 3022 27464
rect 4157 27455 4215 27461
rect 4157 27421 4169 27455
rect 4203 27452 4215 27455
rect 4614 27452 4620 27464
rect 4203 27424 4620 27452
rect 4203 27421 4215 27424
rect 4157 27415 4215 27421
rect 4614 27412 4620 27424
rect 4672 27452 4678 27464
rect 5166 27452 5172 27464
rect 4672 27424 5172 27452
rect 4672 27412 4678 27424
rect 5166 27412 5172 27424
rect 5224 27412 5230 27464
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27285 1639 27319
rect 1581 27279 1639 27285
rect 2130 27276 2136 27328
rect 2188 27316 2194 27328
rect 2498 27316 2504 27328
rect 2188 27288 2504 27316
rect 2188 27276 2194 27288
rect 2498 27276 2504 27288
rect 2556 27276 2562 27328
rect 10134 27316 10140 27328
rect 10095 27288 10140 27316
rect 10134 27276 10140 27288
rect 10192 27276 10198 27328
rect 1104 27226 10856 27248
rect 1104 27174 4213 27226
rect 4265 27174 4277 27226
rect 4329 27174 4341 27226
rect 4393 27174 4405 27226
rect 4457 27174 4469 27226
rect 4521 27174 7477 27226
rect 7529 27174 7541 27226
rect 7593 27174 7605 27226
rect 7657 27174 7669 27226
rect 7721 27174 7733 27226
rect 7785 27174 10856 27226
rect 1104 27152 10856 27174
rect 2961 27115 3019 27121
rect 2961 27112 2973 27115
rect 1872 27084 2973 27112
rect 842 27004 848 27056
rect 900 27044 906 27056
rect 1581 27047 1639 27053
rect 1581 27044 1593 27047
rect 900 27016 1593 27044
rect 900 27004 906 27016
rect 1581 27013 1593 27016
rect 1627 27013 1639 27047
rect 1581 27007 1639 27013
rect 1872 26985 1900 27084
rect 2961 27081 2973 27084
rect 3007 27081 3019 27115
rect 2961 27075 3019 27081
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26945 1915 26979
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 1857 26939 1915 26945
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 3142 26976 3148 26988
rect 3103 26948 3148 26976
rect 3142 26936 3148 26948
rect 3200 26936 3206 26988
rect 1854 26800 1860 26852
rect 1912 26840 1918 26852
rect 2409 26843 2467 26849
rect 2409 26840 2421 26843
rect 1912 26812 2421 26840
rect 1912 26800 1918 26812
rect 2409 26809 2421 26812
rect 2455 26809 2467 26843
rect 2409 26803 2467 26809
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5845 26682
rect 5897 26630 5909 26682
rect 5961 26630 5973 26682
rect 6025 26630 6037 26682
rect 6089 26630 6101 26682
rect 6153 26630 9109 26682
rect 9161 26630 9173 26682
rect 9225 26630 9237 26682
rect 9289 26630 9301 26682
rect 9353 26630 9365 26682
rect 9417 26630 10856 26682
rect 1104 26608 10856 26630
rect 1486 26568 1492 26580
rect 1447 26540 1492 26568
rect 1486 26528 1492 26540
rect 1544 26528 1550 26580
rect 2498 26528 2504 26580
rect 2556 26568 2562 26580
rect 2869 26571 2927 26577
rect 2869 26568 2881 26571
rect 2556 26540 2881 26568
rect 2556 26528 2562 26540
rect 2869 26537 2881 26540
rect 2915 26537 2927 26571
rect 2869 26531 2927 26537
rect 566 26460 572 26512
rect 624 26500 630 26512
rect 2133 26503 2191 26509
rect 2133 26500 2145 26503
rect 624 26472 2145 26500
rect 624 26460 630 26472
rect 2133 26469 2145 26472
rect 2179 26469 2191 26503
rect 2133 26463 2191 26469
rect 2682 26432 2688 26444
rect 1688 26404 2688 26432
rect 1688 26373 1716 26404
rect 2682 26392 2688 26404
rect 2740 26392 2746 26444
rect 10134 26432 10140 26444
rect 10095 26404 10140 26432
rect 10134 26392 10140 26404
rect 10192 26392 10198 26444
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26333 1731 26367
rect 1673 26327 1731 26333
rect 1762 26324 1768 26376
rect 1820 26324 1826 26376
rect 2222 26364 2228 26376
rect 2183 26336 2228 26364
rect 2222 26324 2228 26336
rect 2280 26324 2286 26376
rect 3050 26364 3056 26376
rect 3011 26336 3056 26364
rect 3050 26324 3056 26336
rect 3108 26324 3114 26376
rect 1780 26296 1808 26324
rect 3326 26296 3332 26308
rect 1780 26268 3332 26296
rect 3326 26256 3332 26268
rect 3384 26256 3390 26308
rect 1104 26138 10856 26160
rect 1104 26086 4213 26138
rect 4265 26086 4277 26138
rect 4329 26086 4341 26138
rect 4393 26086 4405 26138
rect 4457 26086 4469 26138
rect 4521 26086 7477 26138
rect 7529 26086 7541 26138
rect 7593 26086 7605 26138
rect 7657 26086 7669 26138
rect 7721 26086 7733 26138
rect 7785 26086 10856 26138
rect 1104 26064 10856 26086
rect 2222 26024 2228 26036
rect 2183 25996 2228 26024
rect 2222 25984 2228 25996
rect 2280 25984 2286 26036
rect 2682 26024 2688 26036
rect 2643 25996 2688 26024
rect 2682 25984 2688 25996
rect 2740 25984 2746 26036
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 1486 25848 1492 25900
rect 1544 25888 1550 25900
rect 2041 25891 2099 25897
rect 2041 25888 2053 25891
rect 1544 25860 2053 25888
rect 1544 25848 1550 25860
rect 2041 25857 2053 25860
rect 2087 25857 2099 25891
rect 2866 25888 2872 25900
rect 2827 25860 2872 25888
rect 2041 25851 2099 25857
rect 2866 25848 2872 25860
rect 2924 25848 2930 25900
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 2130 25684 2136 25696
rect 1627 25656 2136 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 2130 25644 2136 25656
rect 2188 25644 2194 25696
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5845 25594
rect 5897 25542 5909 25594
rect 5961 25542 5973 25594
rect 6025 25542 6037 25594
rect 6089 25542 6101 25594
rect 6153 25542 9109 25594
rect 9161 25542 9173 25594
rect 9225 25542 9237 25594
rect 9289 25542 9301 25594
rect 9353 25542 9365 25594
rect 9417 25542 10856 25594
rect 1104 25520 10856 25542
rect 1949 25483 2007 25489
rect 1949 25449 1961 25483
rect 1995 25480 2007 25483
rect 3694 25480 3700 25492
rect 1995 25452 3700 25480
rect 1995 25449 2007 25452
rect 1949 25443 2007 25449
rect 3694 25440 3700 25452
rect 3752 25440 3758 25492
rect 10134 25480 10140 25492
rect 10095 25452 10140 25480
rect 10134 25440 10140 25452
rect 10192 25440 10198 25492
rect 1949 25279 2007 25285
rect 1949 25245 1961 25279
rect 1995 25276 2007 25279
rect 2593 25279 2651 25285
rect 1995 25248 2452 25276
rect 1995 25245 2007 25248
rect 1949 25239 2007 25245
rect 2424 25149 2452 25248
rect 2593 25245 2605 25279
rect 2639 25276 2651 25279
rect 2774 25276 2780 25288
rect 2639 25248 2780 25276
rect 2639 25245 2651 25248
rect 2593 25239 2651 25245
rect 2774 25236 2780 25248
rect 2832 25236 2838 25288
rect 2409 25143 2467 25149
rect 2409 25109 2421 25143
rect 2455 25109 2467 25143
rect 2409 25103 2467 25109
rect 1104 25050 10856 25072
rect 1104 24998 4213 25050
rect 4265 24998 4277 25050
rect 4329 24998 4341 25050
rect 4393 24998 4405 25050
rect 4457 24998 4469 25050
rect 4521 24998 7477 25050
rect 7529 24998 7541 25050
rect 7593 24998 7605 25050
rect 7657 24998 7669 25050
rect 7721 24998 7733 25050
rect 7785 24998 10856 25050
rect 1104 24976 10856 24998
rect 1397 24803 1455 24809
rect 1397 24769 1409 24803
rect 1443 24800 1455 24803
rect 1486 24800 1492 24812
rect 1443 24772 1492 24800
rect 1443 24769 1455 24772
rect 1397 24763 1455 24769
rect 1486 24760 1492 24772
rect 1544 24760 1550 24812
rect 2130 24800 2136 24812
rect 2091 24772 2136 24800
rect 2130 24760 2136 24772
rect 2188 24760 2194 24812
rect 2958 24800 2964 24812
rect 2919 24772 2964 24800
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 10134 24800 10140 24812
rect 10095 24772 10140 24800
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 1946 24692 1952 24744
rect 2004 24732 2010 24744
rect 2225 24735 2283 24741
rect 2225 24732 2237 24735
rect 2004 24704 2237 24732
rect 2004 24692 2010 24704
rect 2225 24701 2237 24704
rect 2271 24701 2283 24735
rect 2225 24695 2283 24701
rect 2777 24667 2835 24673
rect 2777 24633 2789 24667
rect 2823 24664 2835 24667
rect 3234 24664 3240 24676
rect 2823 24636 3240 24664
rect 2823 24633 2835 24636
rect 2777 24627 2835 24633
rect 3234 24624 3240 24636
rect 3292 24624 3298 24676
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24596 1639 24599
rect 3418 24596 3424 24608
rect 1627 24568 3424 24596
rect 1627 24565 1639 24568
rect 1581 24559 1639 24565
rect 3418 24556 3424 24568
rect 3476 24556 3482 24608
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5845 24506
rect 5897 24454 5909 24506
rect 5961 24454 5973 24506
rect 6025 24454 6037 24506
rect 6089 24454 6101 24506
rect 6153 24454 9109 24506
rect 9161 24454 9173 24506
rect 9225 24454 9237 24506
rect 9289 24454 9301 24506
rect 9353 24454 9365 24506
rect 9417 24454 10856 24506
rect 1104 24432 10856 24454
rect 1210 24352 1216 24404
rect 1268 24392 1274 24404
rect 1673 24395 1731 24401
rect 1673 24392 1685 24395
rect 1268 24364 1685 24392
rect 1268 24352 1274 24364
rect 1673 24361 1685 24364
rect 1719 24361 1731 24395
rect 1673 24355 1731 24361
rect 2869 24395 2927 24401
rect 2869 24361 2881 24395
rect 2915 24392 2927 24395
rect 11057 24395 11115 24401
rect 11057 24392 11069 24395
rect 2915 24364 11069 24392
rect 2915 24361 2927 24364
rect 2869 24355 2927 24361
rect 11057 24361 11069 24364
rect 11103 24361 11115 24395
rect 11057 24355 11115 24361
rect 3970 24284 3976 24336
rect 4028 24284 4034 24336
rect 1670 24216 1676 24268
rect 1728 24256 1734 24268
rect 3418 24256 3424 24268
rect 1728 24228 2728 24256
rect 1728 24216 1734 24228
rect 2700 24197 2728 24228
rect 2884 24228 3424 24256
rect 2884 24197 2912 24228
rect 3418 24216 3424 24228
rect 3476 24256 3482 24268
rect 3988 24256 4016 24284
rect 3476 24228 4016 24256
rect 3476 24216 3482 24228
rect 1857 24191 1915 24197
rect 1857 24157 1869 24191
rect 1903 24157 1915 24191
rect 1857 24151 1915 24157
rect 2685 24191 2743 24197
rect 2685 24157 2697 24191
rect 2731 24157 2743 24191
rect 2685 24151 2743 24157
rect 2869 24191 2927 24197
rect 2869 24157 2881 24191
rect 2915 24157 2927 24191
rect 3970 24188 3976 24200
rect 3931 24160 3976 24188
rect 2869 24151 2927 24157
rect 1872 24052 1900 24151
rect 3970 24148 3976 24160
rect 4028 24148 4034 24200
rect 2314 24080 2320 24132
rect 2372 24120 2378 24132
rect 2498 24120 2504 24132
rect 2372 24092 2504 24120
rect 2372 24080 2378 24092
rect 2498 24080 2504 24092
rect 2556 24080 2562 24132
rect 2746 24092 3832 24120
rect 2746 24052 2774 24092
rect 1872 24024 2774 24052
rect 3234 24012 3240 24064
rect 3292 24052 3298 24064
rect 3694 24052 3700 24064
rect 3292 24024 3700 24052
rect 3292 24012 3298 24024
rect 3694 24012 3700 24024
rect 3752 24012 3758 24064
rect 3804 24061 3832 24092
rect 3789 24055 3847 24061
rect 3789 24021 3801 24055
rect 3835 24021 3847 24055
rect 3789 24015 3847 24021
rect 1104 23962 10856 23984
rect 1104 23910 4213 23962
rect 4265 23910 4277 23962
rect 4329 23910 4341 23962
rect 4393 23910 4405 23962
rect 4457 23910 4469 23962
rect 4521 23910 7477 23962
rect 7529 23910 7541 23962
rect 7593 23910 7605 23962
rect 7657 23910 7669 23962
rect 7721 23910 7733 23962
rect 7785 23910 10856 23962
rect 1104 23888 10856 23910
rect 3789 23851 3847 23857
rect 2056 23820 3464 23848
rect 1210 23672 1216 23724
rect 1268 23712 1274 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 1268 23684 1409 23712
rect 1268 23672 1274 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 1946 23672 1952 23724
rect 2004 23712 2010 23724
rect 2056 23721 2084 23820
rect 2406 23780 2412 23792
rect 2332 23752 2412 23780
rect 2332 23721 2360 23752
rect 2406 23740 2412 23752
rect 2464 23740 2470 23792
rect 2041 23715 2099 23721
rect 2041 23712 2053 23715
rect 2004 23684 2053 23712
rect 2004 23672 2010 23684
rect 2041 23681 2053 23684
rect 2087 23681 2099 23715
rect 2041 23675 2099 23681
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23681 2375 23715
rect 2317 23675 2375 23681
rect 2498 23672 2504 23724
rect 2556 23712 2562 23724
rect 2961 23715 3019 23721
rect 2961 23712 2973 23715
rect 2556 23684 2973 23712
rect 2556 23672 2562 23684
rect 2961 23681 2973 23684
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 3234 23672 3240 23724
rect 3292 23712 3298 23724
rect 3436 23712 3464 23820
rect 3789 23817 3801 23851
rect 3835 23848 3847 23851
rect 11241 23851 11299 23857
rect 11241 23848 11253 23851
rect 3835 23820 11253 23848
rect 3835 23817 3847 23820
rect 3789 23811 3847 23817
rect 11241 23817 11253 23820
rect 11287 23817 11299 23851
rect 11241 23811 11299 23817
rect 3697 23715 3755 23721
rect 3697 23712 3709 23715
rect 3292 23684 3337 23712
rect 3436 23684 3709 23712
rect 3292 23672 3298 23684
rect 3697 23681 3709 23684
rect 3743 23681 3755 23715
rect 3697 23675 3755 23681
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23681 3939 23715
rect 9858 23712 9864 23724
rect 9819 23684 9864 23712
rect 3881 23675 3939 23681
rect 2409 23647 2467 23653
rect 2409 23613 2421 23647
rect 2455 23644 2467 23647
rect 2455 23616 3372 23644
rect 2455 23613 2467 23616
rect 2409 23607 2467 23613
rect 2961 23579 3019 23585
rect 2961 23545 2973 23579
rect 3007 23545 3019 23579
rect 3344 23576 3372 23616
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3896 23644 3924 23675
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 3476 23616 3924 23644
rect 3476 23604 3482 23616
rect 7374 23576 7380 23588
rect 3344 23548 7380 23576
rect 2961 23539 3019 23545
rect 1394 23468 1400 23520
rect 1452 23508 1458 23520
rect 1581 23511 1639 23517
rect 1581 23508 1593 23511
rect 1452 23480 1593 23508
rect 1452 23468 1458 23480
rect 1581 23477 1593 23480
rect 1627 23477 1639 23511
rect 2976 23508 3004 23539
rect 7374 23536 7380 23548
rect 7432 23536 7438 23588
rect 8938 23508 8944 23520
rect 2976 23480 8944 23508
rect 1581 23471 1639 23477
rect 8938 23468 8944 23480
rect 8996 23468 9002 23520
rect 10042 23508 10048 23520
rect 10003 23480 10048 23508
rect 10042 23468 10048 23480
rect 10100 23468 10106 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5845 23418
rect 5897 23366 5909 23418
rect 5961 23366 5973 23418
rect 6025 23366 6037 23418
rect 6089 23366 6101 23418
rect 6153 23366 9109 23418
rect 9161 23366 9173 23418
rect 9225 23366 9237 23418
rect 9289 23366 9301 23418
rect 9353 23366 9365 23418
rect 9417 23366 10856 23418
rect 1104 23344 10856 23366
rect 937 23307 995 23313
rect 937 23273 949 23307
rect 983 23304 995 23307
rect 3878 23304 3884 23316
rect 983 23276 3884 23304
rect 983 23273 995 23276
rect 937 23267 995 23273
rect 3878 23264 3884 23276
rect 3936 23264 3942 23316
rect 9493 23307 9551 23313
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 9858 23304 9864 23316
rect 9539 23276 9864 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 10134 23304 10140 23316
rect 10095 23276 10140 23304
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 1949 23239 2007 23245
rect 1949 23205 1961 23239
rect 1995 23236 2007 23239
rect 2866 23236 2872 23248
rect 1995 23208 2872 23236
rect 1995 23205 2007 23208
rect 1949 23199 2007 23205
rect 2866 23196 2872 23208
rect 2924 23196 2930 23248
rect 3418 23196 3424 23248
rect 3476 23236 3482 23248
rect 3973 23239 4031 23245
rect 3476 23208 3924 23236
rect 3476 23196 3482 23208
rect 2682 23128 2688 23180
rect 2740 23168 2746 23180
rect 2740 23140 3832 23168
rect 2740 23128 2746 23140
rect 1670 23100 1676 23112
rect 1631 23072 1676 23100
rect 1670 23060 1676 23072
rect 1728 23060 1734 23112
rect 1949 23103 2007 23109
rect 1949 23069 1961 23103
rect 1995 23100 2007 23103
rect 2406 23100 2412 23112
rect 1995 23072 2412 23100
rect 1995 23069 2007 23072
rect 1949 23063 2007 23069
rect 2406 23060 2412 23072
rect 2464 23060 2470 23112
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23100 2835 23103
rect 2958 23100 2964 23112
rect 2823 23072 2964 23100
rect 2823 23069 2835 23072
rect 2777 23063 2835 23069
rect 2958 23060 2964 23072
rect 3016 23060 3022 23112
rect 3804 23109 3832 23140
rect 3789 23103 3847 23109
rect 3789 23069 3801 23103
rect 3835 23069 3847 23103
rect 3896 23100 3924 23208
rect 3973 23205 3985 23239
rect 4019 23236 4031 23239
rect 10965 23239 11023 23245
rect 10965 23236 10977 23239
rect 4019 23208 10977 23236
rect 4019 23205 4031 23208
rect 3973 23199 4031 23205
rect 10965 23205 10977 23208
rect 11011 23205 11023 23239
rect 10965 23199 11023 23205
rect 3973 23103 4031 23109
rect 3973 23100 3985 23103
rect 3896 23072 3985 23100
rect 3789 23063 3847 23069
rect 3973 23069 3985 23072
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 9309 23103 9367 23109
rect 9309 23069 9321 23103
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 3053 23035 3111 23041
rect 3053 23001 3065 23035
rect 3099 23001 3111 23035
rect 3053 22995 3111 23001
rect 3068 22964 3096 22995
rect 3234 22992 3240 23044
rect 3292 23032 3298 23044
rect 9324 23032 9352 23063
rect 3292 23004 9352 23032
rect 3292 22992 3298 23004
rect 4614 22964 4620 22976
rect 3068 22936 4620 22964
rect 4614 22924 4620 22936
rect 4672 22924 4678 22976
rect 1104 22874 10856 22896
rect 1104 22822 4213 22874
rect 4265 22822 4277 22874
rect 4329 22822 4341 22874
rect 4393 22822 4405 22874
rect 4457 22822 4469 22874
rect 4521 22822 7477 22874
rect 7529 22822 7541 22874
rect 7593 22822 7605 22874
rect 7657 22822 7669 22874
rect 7721 22822 7733 22874
rect 7785 22822 10856 22874
rect 1104 22800 10856 22822
rect 1489 22763 1547 22769
rect 1489 22729 1501 22763
rect 1535 22760 1547 22763
rect 2222 22760 2228 22772
rect 1535 22732 2228 22760
rect 1535 22729 1547 22732
rect 1489 22723 1547 22729
rect 2222 22720 2228 22732
rect 2280 22720 2286 22772
rect 2498 22760 2504 22772
rect 2424 22732 2504 22760
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22584 1458 22636
rect 2130 22584 2136 22636
rect 2188 22624 2194 22636
rect 2424 22633 2452 22732
rect 2498 22720 2504 22732
rect 2556 22720 2562 22772
rect 3050 22720 3056 22772
rect 3108 22760 3114 22772
rect 3418 22760 3424 22772
rect 3108 22732 3424 22760
rect 3108 22720 3114 22732
rect 3418 22720 3424 22732
rect 3476 22720 3482 22772
rect 3510 22720 3516 22772
rect 3568 22760 3574 22772
rect 3881 22763 3939 22769
rect 3881 22760 3893 22763
rect 3568 22732 3893 22760
rect 3568 22720 3574 22732
rect 3881 22729 3893 22732
rect 3927 22729 3939 22763
rect 3881 22723 3939 22729
rect 2866 22652 2872 22704
rect 2924 22692 2930 22704
rect 6270 22692 6276 22704
rect 2924 22664 6276 22692
rect 2924 22652 2930 22664
rect 6270 22652 6276 22664
rect 6328 22652 6334 22704
rect 2409 22627 2467 22633
rect 2409 22624 2421 22627
rect 2188 22596 2421 22624
rect 2188 22584 2194 22596
rect 2409 22593 2421 22596
rect 2455 22593 2467 22627
rect 2409 22587 2467 22593
rect 3418 22584 3424 22636
rect 3476 22624 3482 22636
rect 4065 22627 4123 22633
rect 4065 22624 4077 22627
rect 3476 22596 4077 22624
rect 3476 22584 3482 22596
rect 4065 22593 4077 22596
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 9766 22584 9772 22636
rect 9824 22624 9830 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9824 22596 9873 22624
rect 9824 22584 9830 22596
rect 9861 22593 9873 22596
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 2498 22516 2504 22568
rect 2556 22556 2562 22568
rect 2777 22559 2835 22565
rect 2777 22556 2789 22559
rect 2556 22528 2789 22556
rect 2556 22516 2562 22528
rect 2777 22525 2789 22528
rect 2823 22525 2835 22559
rect 2777 22519 2835 22525
rect 2406 22448 2412 22500
rect 2464 22488 2470 22500
rect 2682 22488 2688 22500
rect 2464 22460 2688 22488
rect 2464 22448 2470 22460
rect 2682 22448 2688 22460
rect 2740 22448 2746 22500
rect 10042 22488 10048 22500
rect 10003 22460 10048 22488
rect 10042 22448 10048 22460
rect 10100 22448 10106 22500
rect 1104 22330 10856 22352
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5845 22330
rect 5897 22278 5909 22330
rect 5961 22278 5973 22330
rect 6025 22278 6037 22330
rect 6089 22278 6101 22330
rect 6153 22278 9109 22330
rect 9161 22278 9173 22330
rect 9225 22278 9237 22330
rect 9289 22278 9301 22330
rect 9353 22278 9365 22330
rect 9417 22278 10856 22330
rect 1104 22256 10856 22278
rect 2961 22219 3019 22225
rect 2961 22216 2973 22219
rect 2884 22188 2973 22216
rect 2884 22094 2912 22188
rect 2961 22185 2973 22188
rect 3007 22185 3019 22219
rect 2961 22179 3019 22185
rect 3050 22176 3056 22228
rect 3108 22216 3114 22228
rect 3786 22216 3792 22228
rect 3108 22188 3792 22216
rect 3108 22176 3114 22188
rect 3786 22176 3792 22188
rect 3844 22176 3850 22228
rect 1118 22040 1124 22092
rect 1176 22080 1182 22092
rect 1581 22083 1639 22089
rect 1581 22080 1593 22083
rect 1176 22052 1593 22080
rect 1176 22040 1182 22052
rect 1581 22049 1593 22052
rect 1627 22049 1639 22083
rect 2884 22080 3004 22094
rect 1581 22043 1639 22049
rect 1688 22052 3004 22080
rect 1688 22021 1716 22052
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 21981 1731 22015
rect 2314 22012 2320 22024
rect 2275 21984 2320 22012
rect 1673 21975 1731 21981
rect 2314 21972 2320 21984
rect 2372 21972 2378 22024
rect 2406 21972 2412 22024
rect 2464 22012 2470 22024
rect 3142 22012 3148 22024
rect 2464 21984 2509 22012
rect 3103 21984 3148 22012
rect 2464 21972 2470 21984
rect 3142 21972 3148 21984
rect 3200 21972 3206 22024
rect 9217 22015 9275 22021
rect 9217 22012 9229 22015
rect 6886 21984 9229 22012
rect 2746 21916 4752 21944
rect 2409 21879 2467 21885
rect 2409 21845 2421 21879
rect 2455 21876 2467 21879
rect 2746 21876 2774 21916
rect 2455 21848 2774 21876
rect 4724 21876 4752 21916
rect 4798 21904 4804 21956
rect 4856 21944 4862 21956
rect 6886 21944 6914 21984
rect 9217 21981 9229 21984
rect 9263 21981 9275 22015
rect 9858 22012 9864 22024
rect 9819 21984 9864 22012
rect 9217 21975 9275 21981
rect 9858 21972 9864 21984
rect 9916 21972 9922 22024
rect 4856 21916 6914 21944
rect 4856 21904 4862 21916
rect 7282 21876 7288 21888
rect 4724 21848 7288 21876
rect 2455 21845 2467 21848
rect 2409 21839 2467 21845
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 9401 21879 9459 21885
rect 9401 21845 9413 21879
rect 9447 21876 9459 21879
rect 9766 21876 9772 21888
rect 9447 21848 9772 21876
rect 9447 21845 9459 21848
rect 9401 21839 9459 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 1104 21786 10856 21808
rect 1104 21734 4213 21786
rect 4265 21734 4277 21786
rect 4329 21734 4341 21786
rect 4393 21734 4405 21786
rect 4457 21734 4469 21786
rect 4521 21734 7477 21786
rect 7529 21734 7541 21786
rect 7593 21734 7605 21786
rect 7657 21734 7669 21786
rect 7721 21734 7733 21786
rect 7785 21734 10856 21786
rect 1104 21712 10856 21734
rect 2958 21672 2964 21684
rect 2919 21644 2964 21672
rect 2958 21632 2964 21644
rect 3016 21632 3022 21684
rect 1486 21564 1492 21616
rect 1544 21604 1550 21616
rect 4798 21604 4804 21616
rect 1544 21576 4804 21604
rect 1544 21564 1550 21576
rect 4798 21564 4804 21576
rect 4856 21564 4862 21616
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21496 1458 21548
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 3050 21536 3056 21548
rect 2547 21508 3056 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 3050 21496 3056 21508
rect 3108 21496 3114 21548
rect 9766 21496 9772 21548
rect 9824 21536 9830 21548
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 9824 21508 9873 21536
rect 9824 21496 9830 21508
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 9861 21499 9919 21505
rect 2222 21360 2228 21412
rect 2280 21400 2286 21412
rect 2280 21372 2636 21400
rect 2280 21360 2286 21372
rect 1581 21335 1639 21341
rect 1581 21301 1593 21335
rect 1627 21332 1639 21335
rect 2498 21332 2504 21344
rect 1627 21304 2504 21332
rect 1627 21301 1639 21304
rect 1581 21295 1639 21301
rect 2498 21292 2504 21304
rect 2556 21292 2562 21344
rect 2608 21341 2636 21372
rect 2593 21335 2651 21341
rect 2593 21301 2605 21335
rect 2639 21301 2651 21335
rect 10042 21332 10048 21344
rect 10003 21304 10048 21332
rect 2593 21295 2651 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5845 21242
rect 5897 21190 5909 21242
rect 5961 21190 5973 21242
rect 6025 21190 6037 21242
rect 6089 21190 6101 21242
rect 6153 21190 9109 21242
rect 9161 21190 9173 21242
rect 9225 21190 9237 21242
rect 9289 21190 9301 21242
rect 9353 21190 9365 21242
rect 9417 21190 10856 21242
rect 1104 21168 10856 21190
rect 1026 21088 1032 21140
rect 1084 21128 1090 21140
rect 2225 21131 2283 21137
rect 2225 21128 2237 21131
rect 1084 21100 2237 21128
rect 1084 21088 1090 21100
rect 2225 21097 2237 21100
rect 2271 21097 2283 21131
rect 2225 21091 2283 21097
rect 3053 21131 3111 21137
rect 3053 21097 3065 21131
rect 3099 21128 3111 21131
rect 3694 21128 3700 21140
rect 3099 21100 3700 21128
rect 3099 21097 3111 21100
rect 3053 21091 3111 21097
rect 3694 21088 3700 21100
rect 3752 21088 3758 21140
rect 4062 21088 4068 21140
rect 4120 21088 4126 21140
rect 9858 21128 9864 21140
rect 9819 21100 9864 21128
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 3789 21063 3847 21069
rect 3789 21029 3801 21063
rect 3835 21029 3847 21063
rect 3789 21023 3847 21029
rect 3804 20992 3832 21023
rect 2424 20964 3832 20992
rect 2424 20933 2452 20964
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 2409 20927 2467 20933
rect 1719 20896 2360 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 2332 20856 2360 20896
rect 2409 20893 2421 20927
rect 2455 20893 2467 20927
rect 2409 20887 2467 20893
rect 2498 20884 2504 20936
rect 2556 20924 2562 20936
rect 2869 20927 2927 20933
rect 2869 20924 2881 20927
rect 2556 20896 2881 20924
rect 2556 20884 2562 20896
rect 2869 20893 2881 20896
rect 2915 20893 2927 20927
rect 3970 20924 3976 20936
rect 3931 20896 3976 20924
rect 2869 20887 2927 20893
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 3142 20856 3148 20868
rect 2332 20828 3148 20856
rect 3142 20816 3148 20828
rect 3200 20816 3206 20868
rect 3786 20816 3792 20868
rect 3844 20856 3850 20868
rect 4080 20856 4108 21088
rect 10045 20927 10103 20933
rect 10045 20893 10057 20927
rect 10091 20924 10103 20927
rect 11149 20927 11207 20933
rect 11149 20924 11161 20927
rect 10091 20896 11161 20924
rect 10091 20893 10103 20896
rect 10045 20887 10103 20893
rect 11149 20893 11161 20896
rect 11195 20893 11207 20927
rect 11149 20887 11207 20893
rect 3844 20828 4108 20856
rect 3844 20816 3850 20828
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20788 1639 20791
rect 4062 20788 4068 20800
rect 1627 20760 4068 20788
rect 1627 20757 1639 20760
rect 1581 20751 1639 20757
rect 4062 20748 4068 20760
rect 4120 20748 4126 20800
rect 1104 20698 10856 20720
rect 1104 20646 4213 20698
rect 4265 20646 4277 20698
rect 4329 20646 4341 20698
rect 4393 20646 4405 20698
rect 4457 20646 4469 20698
rect 4521 20646 7477 20698
rect 7529 20646 7541 20698
rect 7593 20646 7605 20698
rect 7657 20646 7669 20698
rect 7721 20646 7733 20698
rect 7785 20646 10856 20698
rect 1104 20624 10856 20646
rect 3142 20584 3148 20596
rect 3103 20556 3148 20584
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20448 2099 20451
rect 2685 20451 2743 20457
rect 2087 20420 2544 20448
rect 2087 20417 2099 20420
rect 2041 20411 2099 20417
rect 2516 20321 2544 20420
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2685 20411 2743 20417
rect 2700 20380 2728 20411
rect 2774 20408 2780 20460
rect 2832 20448 2838 20460
rect 3329 20451 3387 20457
rect 3329 20448 3341 20451
rect 2832 20420 3341 20448
rect 2832 20408 2838 20420
rect 3329 20417 3341 20420
rect 3375 20417 3387 20451
rect 3329 20411 3387 20417
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 9861 20451 9919 20457
rect 9861 20448 9873 20451
rect 9732 20420 9873 20448
rect 9732 20408 9738 20420
rect 9861 20417 9873 20420
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 2958 20380 2964 20392
rect 2700 20352 2964 20380
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 2501 20315 2559 20321
rect 2501 20281 2513 20315
rect 2547 20281 2559 20315
rect 3418 20312 3424 20324
rect 2501 20275 2559 20281
rect 2746 20284 3424 20312
rect 1949 20247 2007 20253
rect 1949 20213 1961 20247
rect 1995 20244 2007 20247
rect 2746 20244 2774 20284
rect 3418 20272 3424 20284
rect 3476 20272 3482 20324
rect 10042 20312 10048 20324
rect 10003 20284 10048 20312
rect 10042 20272 10048 20284
rect 10100 20272 10106 20324
rect 1995 20216 2774 20244
rect 1995 20213 2007 20216
rect 1949 20207 2007 20213
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5845 20154
rect 5897 20102 5909 20154
rect 5961 20102 5973 20154
rect 6025 20102 6037 20154
rect 6089 20102 6101 20154
rect 6153 20102 9109 20154
rect 9161 20102 9173 20154
rect 9225 20102 9237 20154
rect 9289 20102 9301 20154
rect 9353 20102 9365 20154
rect 9417 20102 10856 20154
rect 1104 20080 10856 20102
rect 1857 20043 1915 20049
rect 1857 20009 1869 20043
rect 1903 20040 1915 20043
rect 3786 20040 3792 20052
rect 1903 20012 3792 20040
rect 1903 20009 1915 20012
rect 1857 20003 1915 20009
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 1857 19839 1915 19845
rect 1857 19805 1869 19839
rect 1903 19805 1915 19839
rect 1857 19799 1915 19805
rect 2501 19839 2559 19845
rect 2501 19805 2513 19839
rect 2547 19836 2559 19839
rect 2774 19836 2780 19848
rect 2547 19808 2780 19836
rect 2547 19805 2559 19808
rect 2501 19799 2559 19805
rect 1872 19768 1900 19799
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 3142 19836 3148 19848
rect 3103 19808 3148 19836
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 9858 19836 9864 19848
rect 9819 19808 9864 19836
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 1872 19740 3004 19768
rect 1854 19660 1860 19712
rect 1912 19700 1918 19712
rect 2976 19709 3004 19740
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 1912 19672 2329 19700
rect 1912 19660 1918 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 2317 19663 2375 19669
rect 2961 19703 3019 19709
rect 2961 19669 2973 19703
rect 3007 19669 3019 19703
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 2961 19663 3019 19669
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 1104 19610 10856 19632
rect 1104 19558 4213 19610
rect 4265 19558 4277 19610
rect 4329 19558 4341 19610
rect 4393 19558 4405 19610
rect 4457 19558 4469 19610
rect 4521 19558 7477 19610
rect 7529 19558 7541 19610
rect 7593 19558 7605 19610
rect 7657 19558 7669 19610
rect 7721 19558 7733 19610
rect 7785 19558 10856 19610
rect 1104 19536 10856 19558
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 9861 19499 9919 19505
rect 9861 19496 9873 19499
rect 9824 19468 9873 19496
rect 9824 19456 9830 19468
rect 9861 19465 9873 19468
rect 9907 19465 9919 19499
rect 9861 19459 9919 19465
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 2317 19363 2375 19369
rect 2317 19329 2329 19363
rect 2363 19360 2375 19363
rect 2958 19360 2964 19372
rect 2363 19332 2964 19360
rect 2363 19329 2375 19332
rect 2317 19323 2375 19329
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19360 10103 19363
rect 11057 19363 11115 19369
rect 11057 19360 11069 19363
rect 10091 19332 11069 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 11057 19329 11069 19332
rect 11103 19329 11115 19363
rect 11057 19323 11115 19329
rect 1857 19227 1915 19233
rect 1857 19193 1869 19227
rect 1903 19224 1915 19227
rect 3602 19224 3608 19236
rect 1903 19196 3608 19224
rect 1903 19193 1915 19196
rect 1857 19187 1915 19193
rect 3602 19184 3608 19196
rect 3660 19184 3666 19236
rect 2498 19156 2504 19168
rect 2459 19128 2504 19156
rect 2498 19116 2504 19128
rect 2556 19116 2562 19168
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5845 19066
rect 5897 19014 5909 19066
rect 5961 19014 5973 19066
rect 6025 19014 6037 19066
rect 6089 19014 6101 19066
rect 6153 19014 9109 19066
rect 9161 19014 9173 19066
rect 9225 19014 9237 19066
rect 9289 19014 9301 19066
rect 9353 19014 9365 19066
rect 9417 19014 10856 19066
rect 1104 18992 10856 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 9858 18952 9864 18964
rect 9447 18924 9864 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 2130 18776 2136 18828
rect 2188 18816 2194 18828
rect 3053 18819 3111 18825
rect 3053 18816 3065 18819
rect 2188 18788 3065 18816
rect 2188 18776 2194 18788
rect 3053 18785 3065 18788
rect 3099 18816 3111 18819
rect 4062 18816 4068 18828
rect 3099 18788 4068 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 2406 18748 2412 18760
rect 2367 18720 2412 18748
rect 1765 18711 1823 18717
rect 1780 18680 1808 18711
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 2682 18708 2688 18760
rect 2740 18748 2746 18760
rect 3970 18748 3976 18760
rect 2740 18720 3188 18748
rect 3931 18720 3976 18748
rect 2740 18708 2746 18720
rect 3160 18680 3188 18720
rect 3970 18708 3976 18720
rect 4028 18708 4034 18760
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 6886 18720 9229 18748
rect 6886 18680 6914 18720
rect 9217 18717 9229 18720
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9766 18708 9772 18760
rect 9824 18748 9830 18760
rect 9861 18751 9919 18757
rect 9861 18748 9873 18751
rect 9824 18720 9873 18748
rect 9824 18708 9830 18720
rect 9861 18717 9873 18720
rect 9907 18717 9919 18751
rect 9861 18711 9919 18717
rect 1780 18652 2774 18680
rect 3160 18652 6914 18680
rect 2746 18612 2774 18652
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 2746 18584 3801 18612
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 10042 18612 10048 18624
rect 10003 18584 10048 18612
rect 3789 18575 3847 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 1104 18522 10856 18544
rect 1104 18470 4213 18522
rect 4265 18470 4277 18522
rect 4329 18470 4341 18522
rect 4393 18470 4405 18522
rect 4457 18470 4469 18522
rect 4521 18470 7477 18522
rect 7529 18470 7541 18522
rect 7593 18470 7605 18522
rect 7657 18470 7669 18522
rect 7721 18470 7733 18522
rect 7785 18470 10856 18522
rect 1104 18448 10856 18470
rect 1670 18408 1676 18420
rect 1631 18380 1676 18408
rect 1670 18368 1676 18380
rect 1728 18368 1734 18420
rect 2406 18408 2412 18420
rect 2367 18380 2412 18408
rect 2406 18368 2412 18380
rect 2464 18368 2470 18420
rect 9401 18411 9459 18417
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 9674 18408 9680 18420
rect 9447 18380 9680 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 2222 18300 2228 18352
rect 2280 18340 2286 18352
rect 2593 18343 2651 18349
rect 2593 18340 2605 18343
rect 2280 18312 2605 18340
rect 2280 18300 2286 18312
rect 2593 18309 2605 18312
rect 2639 18309 2651 18343
rect 2593 18303 2651 18309
rect 2777 18343 2835 18349
rect 2777 18309 2789 18343
rect 2823 18340 2835 18343
rect 3050 18340 3056 18352
rect 2823 18312 3056 18340
rect 2823 18309 2835 18312
rect 2777 18303 2835 18309
rect 3050 18300 3056 18312
rect 3108 18300 3114 18352
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18241 1823 18275
rect 1765 18235 1823 18241
rect 1780 18204 1808 18235
rect 2406 18232 2412 18284
rect 2464 18272 2470 18284
rect 2682 18272 2688 18284
rect 2464 18244 2688 18272
rect 2464 18232 2470 18244
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 3418 18272 3424 18284
rect 3379 18244 3424 18272
rect 3418 18232 3424 18244
rect 3476 18232 3482 18284
rect 9217 18275 9275 18281
rect 9217 18272 9229 18275
rect 6886 18244 9229 18272
rect 3786 18204 3792 18216
rect 1780 18176 3792 18204
rect 3786 18164 3792 18176
rect 3844 18164 3850 18216
rect 1854 18096 1860 18148
rect 1912 18136 1918 18148
rect 6886 18136 6914 18244
rect 9217 18241 9229 18244
rect 9263 18241 9275 18275
rect 9217 18235 9275 18241
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18272 9919 18275
rect 9950 18272 9956 18284
rect 9907 18244 9956 18272
rect 9907 18241 9919 18244
rect 9861 18235 9919 18241
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 1912 18108 6914 18136
rect 1912 18096 1918 18108
rect 3234 18068 3240 18080
rect 3195 18040 3240 18068
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5845 17978
rect 5897 17926 5909 17978
rect 5961 17926 5973 17978
rect 6025 17926 6037 17978
rect 6089 17926 6101 17978
rect 6153 17926 9109 17978
rect 9161 17926 9173 17978
rect 9225 17926 9237 17978
rect 9289 17926 9301 17978
rect 9353 17926 9365 17978
rect 9417 17926 10856 17978
rect 1104 17904 10856 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 3786 17864 3792 17876
rect 3747 17836 3792 17864
rect 3786 17824 3792 17836
rect 3844 17824 3850 17876
rect 1578 17756 1584 17808
rect 1636 17796 1642 17808
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 1636 17768 2605 17796
rect 1636 17756 1642 17768
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 2593 17759 2651 17765
rect 3234 17728 3240 17740
rect 2056 17700 3240 17728
rect 2056 17669 2084 17700
rect 3234 17688 3240 17700
rect 3292 17688 3298 17740
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17629 2099 17663
rect 2498 17660 2504 17672
rect 2459 17632 2504 17660
rect 2041 17623 2099 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 3970 17660 3976 17672
rect 3931 17632 3976 17660
rect 3970 17620 3976 17632
rect 4028 17620 4034 17672
rect 9858 17660 9864 17672
rect 9819 17632 9864 17660
rect 9858 17620 9864 17632
rect 9916 17620 9922 17672
rect 10042 17524 10048 17536
rect 10003 17496 10048 17524
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 1104 17434 10856 17456
rect 1104 17382 4213 17434
rect 4265 17382 4277 17434
rect 4329 17382 4341 17434
rect 4393 17382 4405 17434
rect 4457 17382 4469 17434
rect 4521 17382 7477 17434
rect 7529 17382 7541 17434
rect 7593 17382 7605 17434
rect 7657 17382 7669 17434
rect 7721 17382 7733 17434
rect 7785 17382 10856 17434
rect 1104 17360 10856 17382
rect 9950 17320 9956 17332
rect 9911 17292 9956 17320
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17144 1458 17196
rect 1486 17144 1492 17196
rect 1544 17184 1550 17196
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 1544 17156 2237 17184
rect 1544 17144 1550 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2866 17184 2872 17196
rect 2827 17156 2872 17184
rect 2225 17147 2283 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10183 17156 10977 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1820 16952 2053 16980
rect 1820 16940 1826 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 2222 16940 2228 16992
rect 2280 16980 2286 16992
rect 2685 16983 2743 16989
rect 2685 16980 2697 16983
rect 2280 16952 2697 16980
rect 2280 16940 2286 16952
rect 2685 16949 2697 16952
rect 2731 16949 2743 16983
rect 2685 16943 2743 16949
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5845 16890
rect 5897 16838 5909 16890
rect 5961 16838 5973 16890
rect 6025 16838 6037 16890
rect 6089 16838 6101 16890
rect 6153 16838 9109 16890
rect 9161 16838 9173 16890
rect 9225 16838 9237 16890
rect 9289 16838 9301 16890
rect 9353 16838 9365 16890
rect 9417 16838 10856 16890
rect 1104 16816 10856 16838
rect 2222 16640 2228 16652
rect 2148 16612 2228 16640
rect 2148 16581 2176 16612
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2774 16572 2780 16584
rect 2735 16544 2780 16572
rect 2133 16535 2191 16541
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 9217 16575 9275 16581
rect 9217 16572 9229 16575
rect 6886 16544 9229 16572
rect 2041 16507 2099 16513
rect 2041 16473 2053 16507
rect 2087 16504 2099 16507
rect 2314 16504 2320 16516
rect 2087 16476 2320 16504
rect 2087 16473 2099 16476
rect 2041 16467 2099 16473
rect 2314 16464 2320 16476
rect 2372 16464 2378 16516
rect 2498 16464 2504 16516
rect 2556 16504 2562 16516
rect 6886 16504 6914 16544
rect 9217 16541 9229 16544
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9732 16544 9873 16572
rect 9732 16532 9738 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 2556 16476 6914 16504
rect 2556 16464 2562 16476
rect 2590 16436 2596 16448
rect 2551 16408 2596 16436
rect 2590 16396 2596 16408
rect 2648 16396 2654 16448
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9766 16436 9772 16448
rect 9447 16408 9772 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 1104 16346 10856 16368
rect 1104 16294 4213 16346
rect 4265 16294 4277 16346
rect 4329 16294 4341 16346
rect 4393 16294 4405 16346
rect 4457 16294 4469 16346
rect 4521 16294 7477 16346
rect 7529 16294 7541 16346
rect 7593 16294 7605 16346
rect 7657 16294 7669 16346
rect 7721 16294 7733 16346
rect 7785 16294 10856 16346
rect 1104 16272 10856 16294
rect 1949 16235 2007 16241
rect 1949 16201 1961 16235
rect 1995 16232 2007 16235
rect 2130 16232 2136 16244
rect 1995 16204 2136 16232
rect 1995 16201 2007 16204
rect 1949 16195 2007 16201
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2240 16204 2605 16232
rect 1670 16124 1676 16176
rect 1728 16164 1734 16176
rect 1728 16136 1992 16164
rect 1728 16124 1734 16136
rect 1486 16096 1492 16108
rect 1447 16068 1492 16096
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 1762 16096 1768 16108
rect 1723 16068 1768 16096
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 1964 16096 1992 16136
rect 2240 16096 2268 16204
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 11057 16235 11115 16241
rect 11057 16232 11069 16235
rect 2593 16195 2651 16201
rect 6886 16204 11069 16232
rect 2424 16136 2774 16164
rect 1964 16068 2268 16096
rect 2314 16056 2320 16108
rect 2372 16096 2378 16108
rect 2424 16105 2452 16136
rect 2409 16099 2467 16105
rect 2409 16096 2421 16099
rect 2372 16068 2421 16096
rect 2372 16056 2378 16068
rect 2409 16065 2421 16068
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 2501 16102 2559 16105
rect 2501 16099 2636 16102
rect 2501 16065 2513 16099
rect 2547 16074 2636 16099
rect 2547 16065 2559 16074
rect 2501 16059 2559 16065
rect 1673 16031 1731 16037
rect 1673 15997 1685 16031
rect 1719 15997 1731 16031
rect 1673 15991 1731 15997
rect 1688 15904 1716 15991
rect 2038 15988 2044 16040
rect 2096 16028 2102 16040
rect 2608 16028 2636 16074
rect 2746 16096 2774 16136
rect 6886 16096 6914 16204
rect 11057 16201 11069 16204
rect 11103 16201 11115 16235
rect 11057 16195 11115 16201
rect 2746 16068 6914 16096
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 9907 16068 11069 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 11057 16065 11069 16068
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 2096 16000 2636 16028
rect 2777 16031 2835 16037
rect 2096 15988 2102 16000
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 3234 16028 3240 16040
rect 2823 16000 3240 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 2590 15960 2596 15972
rect 1780 15932 2596 15960
rect 1670 15852 1676 15904
rect 1728 15852 1734 15904
rect 1780 15901 1808 15932
rect 2590 15920 2596 15932
rect 2648 15920 2654 15972
rect 1765 15895 1823 15901
rect 1765 15861 1777 15895
rect 1811 15861 1823 15895
rect 1765 15855 1823 15861
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 2501 15895 2559 15901
rect 2501 15892 2513 15895
rect 2464 15864 2513 15892
rect 2464 15852 2470 15864
rect 2501 15861 2513 15864
rect 2547 15861 2559 15895
rect 10042 15892 10048 15904
rect 10003 15864 10048 15892
rect 2501 15855 2559 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5845 15802
rect 5897 15750 5909 15802
rect 5961 15750 5973 15802
rect 6025 15750 6037 15802
rect 6089 15750 6101 15802
rect 6153 15750 9109 15802
rect 9161 15750 9173 15802
rect 9225 15750 9237 15802
rect 9289 15750 9301 15802
rect 9353 15750 9365 15802
rect 9417 15750 10856 15802
rect 1104 15728 10856 15750
rect 1489 15691 1547 15697
rect 1489 15657 1501 15691
rect 1535 15688 1547 15691
rect 1670 15688 1676 15700
rect 1535 15660 1676 15688
rect 1535 15657 1547 15660
rect 1489 15651 1547 15657
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2096 15660 6914 15688
rect 2096 15648 2102 15660
rect 2685 15623 2743 15629
rect 2685 15589 2697 15623
rect 2731 15589 2743 15623
rect 6886 15620 6914 15660
rect 9858 15648 9864 15700
rect 9916 15688 9922 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9916 15660 9965 15688
rect 9916 15648 9922 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 9953 15651 10011 15657
rect 11149 15623 11207 15629
rect 11149 15620 11161 15623
rect 6886 15592 11161 15620
rect 2685 15583 2743 15589
rect 11149 15589 11161 15592
rect 11195 15589 11207 15623
rect 11149 15583 11207 15589
rect 2700 15552 2728 15583
rect 1412 15524 2728 15552
rect 1412 15493 1440 15524
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15453 1455 15487
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1397 15447 1455 15453
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 10134 15484 10140 15496
rect 10095 15456 10140 15484
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 2498 15416 2504 15428
rect 1596 15388 2504 15416
rect 1596 15360 1624 15388
rect 2498 15376 2504 15388
rect 2556 15376 2562 15428
rect 1578 15308 1584 15360
rect 1636 15308 1642 15360
rect 1762 15308 1768 15360
rect 1820 15348 1826 15360
rect 2041 15351 2099 15357
rect 2041 15348 2053 15351
rect 1820 15320 2053 15348
rect 1820 15308 1826 15320
rect 2041 15317 2053 15320
rect 2087 15317 2099 15351
rect 2041 15311 2099 15317
rect 1104 15258 10856 15280
rect 1104 15206 4213 15258
rect 4265 15206 4277 15258
rect 4329 15206 4341 15258
rect 4393 15206 4405 15258
rect 4457 15206 4469 15258
rect 4521 15206 7477 15258
rect 7529 15206 7541 15258
rect 7593 15206 7605 15258
rect 7657 15206 7669 15258
rect 7721 15206 7733 15258
rect 7785 15206 10856 15258
rect 1104 15184 10856 15206
rect 1394 15104 1400 15156
rect 1452 15144 1458 15156
rect 1857 15147 1915 15153
rect 1857 15144 1869 15147
rect 1452 15116 1869 15144
rect 1452 15104 1458 15116
rect 1857 15113 1869 15116
rect 1903 15144 1915 15147
rect 2130 15144 2136 15156
rect 1903 15116 2136 15144
rect 1903 15113 1915 15116
rect 1857 15107 1915 15113
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3050 15144 3056 15156
rect 3007 15116 3056 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 1578 15036 1584 15088
rect 1636 15076 1642 15088
rect 1765 15079 1823 15085
rect 1765 15076 1777 15079
rect 1636 15048 1777 15076
rect 1636 15036 1642 15048
rect 1765 15045 1777 15048
rect 1811 15045 1823 15079
rect 1765 15039 1823 15045
rect 2240 15048 9674 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 1688 14940 1716 14971
rect 1854 14968 1860 15020
rect 1912 15008 1918 15020
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 1912 14980 2053 15008
rect 1912 14968 1918 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 2240 14940 2268 15048
rect 2501 15011 2559 15017
rect 2501 15008 2513 15011
rect 1688 14912 2268 14940
rect 2332 14980 2513 15008
rect 2148 14884 2176 14912
rect 2130 14832 2136 14884
rect 2188 14832 2194 14884
rect 1949 14807 2007 14813
rect 1949 14773 1961 14807
rect 1995 14804 2007 14807
rect 2332 14804 2360 14980
rect 2501 14977 2513 14980
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 2958 15008 2964 15020
rect 2823 14980 2964 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2958 14968 2964 14980
rect 3016 14968 3022 15020
rect 2406 14900 2412 14952
rect 2464 14940 2470 14952
rect 2593 14943 2651 14949
rect 2593 14940 2605 14943
rect 2464 14912 2605 14940
rect 2464 14900 2470 14912
rect 2593 14909 2605 14912
rect 2639 14909 2651 14943
rect 9646 14940 9674 15048
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 9907 14980 11253 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 11241 14977 11253 14980
rect 11287 14977 11299 15011
rect 11241 14971 11299 14977
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 9646 14912 10977 14940
rect 2593 14903 2651 14909
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 10042 14872 10048 14884
rect 10003 14844 10048 14872
rect 10042 14832 10048 14844
rect 10100 14832 10106 14884
rect 2498 14804 2504 14816
rect 1995 14776 2360 14804
rect 2459 14776 2504 14804
rect 1995 14773 2007 14776
rect 1949 14767 2007 14773
rect 2498 14764 2504 14776
rect 2556 14764 2562 14816
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5845 14714
rect 5897 14662 5909 14714
rect 5961 14662 5973 14714
rect 6025 14662 6037 14714
rect 6089 14662 6101 14714
rect 6153 14662 9109 14714
rect 9161 14662 9173 14714
rect 9225 14662 9237 14714
rect 9289 14662 9301 14714
rect 9353 14662 9365 14714
rect 9417 14662 10856 14714
rect 1104 14640 10856 14662
rect 1397 14603 1455 14609
rect 1397 14569 1409 14603
rect 1443 14600 1455 14603
rect 1486 14600 1492 14612
rect 1443 14572 1492 14600
rect 1443 14569 1455 14572
rect 1397 14563 1455 14569
rect 1486 14560 1492 14572
rect 1544 14560 1550 14612
rect 1857 14603 1915 14609
rect 1857 14569 1869 14603
rect 1903 14600 1915 14603
rect 2317 14603 2375 14609
rect 2317 14600 2329 14603
rect 1903 14572 2329 14600
rect 1903 14569 1915 14572
rect 1857 14563 1915 14569
rect 2317 14569 2329 14572
rect 2363 14569 2375 14603
rect 2317 14563 2375 14569
rect 1670 14532 1676 14544
rect 1504 14504 1676 14532
rect 1504 14476 1532 14504
rect 1670 14492 1676 14504
rect 1728 14492 1734 14544
rect 1486 14424 1492 14476
rect 1544 14424 1550 14476
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 1596 14260 1624 14359
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 2501 14399 2559 14405
rect 2501 14396 2513 14399
rect 1728 14368 2513 14396
rect 1728 14356 1734 14368
rect 2501 14365 2513 14368
rect 2547 14365 2559 14399
rect 3142 14396 3148 14408
rect 3103 14368 3148 14396
rect 2501 14359 2559 14365
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 9907 14368 10977 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 1857 14331 1915 14337
rect 1857 14297 1869 14331
rect 1903 14328 1915 14331
rect 1903 14300 3832 14328
rect 1903 14297 1915 14300
rect 1857 14291 1915 14297
rect 3804 14269 3832 14300
rect 2961 14263 3019 14269
rect 2961 14260 2973 14263
rect 1596 14232 2973 14260
rect 2961 14229 2973 14232
rect 3007 14229 3019 14263
rect 2961 14223 3019 14229
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 3789 14223 3847 14229
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 1104 14170 10856 14192
rect 1104 14118 4213 14170
rect 4265 14118 4277 14170
rect 4329 14118 4341 14170
rect 4393 14118 4405 14170
rect 4457 14118 4469 14170
rect 4521 14118 7477 14170
rect 7529 14118 7541 14170
rect 7593 14118 7605 14170
rect 7657 14118 7669 14170
rect 7721 14118 7733 14170
rect 7785 14118 10856 14170
rect 1104 14096 10856 14118
rect 1486 14016 1492 14068
rect 1544 14056 1550 14068
rect 1949 14059 2007 14065
rect 1949 14056 1961 14059
rect 1544 14028 1961 14056
rect 1544 14016 1550 14028
rect 1949 14025 1961 14028
rect 1995 14025 2007 14059
rect 1949 14019 2007 14025
rect 2869 14059 2927 14065
rect 2869 14025 2881 14059
rect 2915 14056 2927 14059
rect 2958 14056 2964 14068
rect 2915 14028 2964 14056
rect 2915 14025 2927 14028
rect 2869 14019 2927 14025
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9674 14056 9680 14068
rect 9447 14028 9680 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 2372 13960 6914 13988
rect 2372 13948 2378 13960
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2700 13929 2728 13960
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2869 13923 2927 13929
rect 2731 13892 2765 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2869 13889 2881 13923
rect 2915 13889 2927 13923
rect 6886 13920 6914 13960
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 6886 13892 9229 13920
rect 2869 13883 2927 13889
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 9907 13892 11161 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 11149 13889 11161 13892
rect 11195 13889 11207 13923
rect 11149 13883 11207 13889
rect 2884 13852 2912 13883
rect 3142 13852 3148 13864
rect 2884 13824 3148 13852
rect 3142 13812 3148 13824
rect 3200 13852 3206 13864
rect 10134 13852 10140 13864
rect 3200 13824 10140 13852
rect 3200 13812 3206 13824
rect 10134 13812 10140 13824
rect 10192 13812 10198 13864
rect 10042 13716 10048 13728
rect 10003 13688 10048 13716
rect 10042 13676 10048 13688
rect 10100 13676 10106 13728
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5845 13626
rect 5897 13574 5909 13626
rect 5961 13574 5973 13626
rect 6025 13574 6037 13626
rect 6089 13574 6101 13626
rect 6153 13574 9109 13626
rect 9161 13574 9173 13626
rect 9225 13574 9237 13626
rect 9289 13574 9301 13626
rect 9353 13574 9365 13626
rect 9417 13574 10856 13626
rect 1104 13552 10856 13574
rect 2961 13447 3019 13453
rect 2961 13413 2973 13447
rect 3007 13444 3019 13447
rect 3234 13444 3240 13456
rect 3007 13416 3240 13444
rect 3007 13413 3019 13416
rect 2961 13407 3019 13413
rect 3234 13404 3240 13416
rect 3292 13404 3298 13456
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 2038 13376 2044 13388
rect 1719 13348 2044 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 2038 13336 2044 13348
rect 2096 13336 2102 13388
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 1762 13200 1768 13252
rect 1820 13240 1826 13252
rect 2038 13240 2044 13252
rect 1820 13212 2044 13240
rect 1820 13200 1826 13212
rect 2038 13200 2044 13212
rect 2096 13200 2102 13252
rect 2774 13240 2780 13252
rect 2735 13212 2780 13240
rect 2774 13200 2780 13212
rect 2832 13200 2838 13252
rect 1104 13082 10856 13104
rect 1104 13030 4213 13082
rect 4265 13030 4277 13082
rect 4329 13030 4341 13082
rect 4393 13030 4405 13082
rect 4457 13030 4469 13082
rect 4521 13030 7477 13082
rect 7529 13030 7541 13082
rect 7593 13030 7605 13082
rect 7657 13030 7669 13082
rect 7721 13030 7733 13082
rect 7785 13030 10856 13082
rect 1104 13008 10856 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1762 12968 1768 12980
rect 1544 12940 1768 12968
rect 1544 12928 1550 12940
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 2777 12971 2835 12977
rect 2777 12937 2789 12971
rect 2823 12968 2835 12971
rect 7834 12968 7840 12980
rect 2823 12940 7840 12968
rect 2823 12937 2835 12940
rect 2777 12931 2835 12937
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2222 12832 2228 12844
rect 1719 12804 2228 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2222 12792 2228 12804
rect 2280 12792 2286 12844
rect 2961 12835 3019 12841
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3418 12832 3424 12844
rect 3007 12804 3424 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 9824 12804 9873 12832
rect 9824 12792 9830 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 1302 12724 1308 12776
rect 1360 12764 1366 12776
rect 1397 12767 1455 12773
rect 1397 12764 1409 12767
rect 1360 12736 1409 12764
rect 1360 12724 1366 12736
rect 1397 12733 1409 12736
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 10042 12628 10048 12640
rect 10003 12600 10048 12628
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5845 12538
rect 5897 12486 5909 12538
rect 5961 12486 5973 12538
rect 6025 12486 6037 12538
rect 6089 12486 6101 12538
rect 6153 12486 9109 12538
rect 9161 12486 9173 12538
rect 9225 12486 9237 12538
rect 9289 12486 9301 12538
rect 9353 12486 9365 12538
rect 9417 12486 10856 12538
rect 1104 12464 10856 12486
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 7926 12424 7932 12436
rect 2823 12396 7932 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 2038 12288 2044 12300
rect 1719 12260 2044 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 3786 12220 3792 12232
rect 3747 12192 3792 12220
rect 2961 12183 3019 12189
rect 2976 12152 3004 12183
rect 3786 12180 3792 12192
rect 3844 12180 3850 12232
rect 9858 12220 9864 12232
rect 9819 12192 9864 12220
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 3878 12152 3884 12164
rect 2976 12124 3884 12152
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 9766 12084 9772 12096
rect 4019 12056 9772 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 9766 12044 9772 12056
rect 9824 12044 9830 12096
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 1104 11994 10856 12016
rect 1104 11942 4213 11994
rect 4265 11942 4277 11994
rect 4329 11942 4341 11994
rect 4393 11942 4405 11994
rect 4457 11942 4469 11994
rect 4521 11942 7477 11994
rect 7529 11942 7541 11994
rect 7593 11942 7605 11994
rect 7657 11942 7669 11994
rect 7721 11942 7733 11994
rect 7785 11942 10856 11994
rect 1104 11920 10856 11942
rect 2777 11883 2835 11889
rect 2777 11849 2789 11883
rect 2823 11880 2835 11883
rect 7190 11880 7196 11892
rect 2823 11852 7196 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 3234 11772 3240 11824
rect 3292 11812 3298 11824
rect 3292 11784 4108 11812
rect 3292 11772 3298 11784
rect 4080 11756 4108 11784
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1762 11744 1768 11756
rect 1719 11716 1768 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 2961 11747 3019 11753
rect 2961 11744 2973 11747
rect 2280 11716 2973 11744
rect 2280 11704 2286 11716
rect 2961 11713 2973 11716
rect 3007 11713 3019 11747
rect 3418 11744 3424 11756
rect 3379 11716 3424 11744
rect 2961 11707 3019 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 4062 11744 4068 11756
rect 3975 11716 4068 11744
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 1360 11648 1409 11676
rect 1360 11636 1366 11648
rect 1397 11645 1409 11648
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 3602 11540 3608 11552
rect 3563 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 9858 11540 9864 11552
rect 4295 11512 9864 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5845 11450
rect 5897 11398 5909 11450
rect 5961 11398 5973 11450
rect 6025 11398 6037 11450
rect 6089 11398 6101 11450
rect 6153 11398 9109 11450
rect 9161 11398 9173 11450
rect 9225 11398 9237 11450
rect 9289 11398 9301 11450
rect 9353 11398 9365 11450
rect 9417 11398 10856 11450
rect 1104 11376 10856 11398
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 3660 11308 9904 11336
rect 3660 11296 3666 11308
rect 3973 11271 4031 11277
rect 3973 11237 3985 11271
rect 4019 11268 4031 11271
rect 9674 11268 9680 11280
rect 4019 11240 9680 11268
rect 4019 11237 4031 11240
rect 3973 11231 4031 11237
rect 9674 11228 9680 11240
rect 9732 11228 9738 11280
rect 1486 11160 1492 11212
rect 1544 11200 1550 11212
rect 1673 11203 1731 11209
rect 1673 11200 1685 11203
rect 1544 11172 1685 11200
rect 1544 11160 1550 11172
rect 1673 11169 1685 11172
rect 1719 11169 1731 11203
rect 1673 11163 1731 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2685 11135 2743 11141
rect 2685 11132 2697 11135
rect 2280 11104 2697 11132
rect 2280 11092 2286 11104
rect 2685 11101 2697 11104
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11132 3847 11135
rect 3878 11132 3884 11144
rect 3835 11104 3884 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 9876 11141 9904 11308
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 9766 11064 9772 11076
rect 2884 11036 9772 11064
rect 2884 11005 2912 11036
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 2869 10999 2927 11005
rect 2869 10965 2881 10999
rect 2915 10965 2927 10999
rect 2869 10959 2927 10965
rect 1104 10906 10856 10928
rect 1104 10854 4213 10906
rect 4265 10854 4277 10906
rect 4329 10854 4341 10906
rect 4393 10854 4405 10906
rect 4457 10854 4469 10906
rect 4521 10854 7477 10906
rect 7529 10854 7541 10906
rect 7593 10854 7605 10906
rect 7657 10854 7669 10906
rect 7721 10854 7733 10906
rect 7785 10854 10856 10906
rect 1104 10832 10856 10854
rect 3421 10727 3479 10733
rect 3421 10693 3433 10727
rect 3467 10724 3479 10727
rect 9030 10724 9036 10736
rect 3467 10696 9036 10724
rect 3467 10693 3479 10696
rect 3421 10687 3479 10693
rect 9030 10684 9036 10696
rect 9088 10684 9094 10736
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2130 10656 2136 10668
rect 1719 10628 2136 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 2130 10616 2136 10628
rect 2188 10616 2194 10668
rect 2961 10659 3019 10665
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3050 10656 3056 10668
rect 3007 10628 3056 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3050 10616 3056 10628
rect 3108 10616 3114 10668
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10656 3295 10659
rect 3970 10656 3976 10668
rect 3283 10628 3976 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 1360 10560 1409 10588
rect 1360 10548 1366 10560
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 3252 10520 3280 10619
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 9732 10628 9873 10656
rect 9732 10616 9738 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 3016 10492 3280 10520
rect 3016 10480 3022 10492
rect 10042 10452 10048 10464
rect 10003 10424 10048 10452
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5845 10362
rect 5897 10310 5909 10362
rect 5961 10310 5973 10362
rect 6025 10310 6037 10362
rect 6089 10310 6101 10362
rect 6153 10310 9109 10362
rect 9161 10310 9173 10362
rect 9225 10310 9237 10362
rect 9289 10310 9301 10362
rect 9353 10310 9365 10362
rect 9417 10310 10856 10362
rect 1104 10288 10856 10310
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 9999 10220 10977 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10965 10217 10977 10220
rect 11011 10217 11023 10251
rect 10965 10211 11023 10217
rect 9493 10183 9551 10189
rect 9493 10149 9505 10183
rect 9539 10180 9551 10183
rect 11057 10183 11115 10189
rect 11057 10180 11069 10183
rect 9539 10152 11069 10180
rect 9539 10149 9551 10152
rect 9493 10143 9551 10149
rect 11057 10149 11069 10152
rect 11103 10149 11115 10183
rect 11057 10143 11115 10149
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 3142 10112 3148 10124
rect 1719 10084 3148 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 3142 10072 3148 10084
rect 3200 10072 3206 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2685 10047 2743 10053
rect 2685 10044 2697 10047
rect 2188 10016 2697 10044
rect 2188 10004 2194 10016
rect 2685 10013 2697 10016
rect 2731 10013 2743 10047
rect 2685 10007 2743 10013
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 4672 10016 9321 10044
rect 4672 10004 4678 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 9309 10007 9367 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 2869 9911 2927 9917
rect 2869 9877 2881 9911
rect 2915 9908 2927 9911
rect 9858 9908 9864 9920
rect 2915 9880 9864 9908
rect 2915 9877 2927 9880
rect 2869 9871 2927 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 1104 9818 10856 9840
rect 1104 9766 4213 9818
rect 4265 9766 4277 9818
rect 4329 9766 4341 9818
rect 4393 9766 4405 9818
rect 4457 9766 4469 9818
rect 4521 9766 7477 9818
rect 7529 9766 7541 9818
rect 7593 9766 7605 9818
rect 7657 9766 7669 9818
rect 7721 9766 7733 9818
rect 7785 9766 10856 9818
rect 1104 9744 10856 9766
rect 2777 9707 2835 9713
rect 2777 9673 2789 9707
rect 2823 9704 2835 9707
rect 3970 9704 3976 9716
rect 2823 9676 3976 9704
rect 2823 9673 2835 9676
rect 2777 9667 2835 9673
rect 3970 9664 3976 9676
rect 4028 9704 4034 9716
rect 10134 9704 10140 9716
rect 4028 9676 10140 9704
rect 4028 9664 4034 9676
rect 10134 9664 10140 9676
rect 10192 9664 10198 9716
rect 2888 9639 2946 9645
rect 2888 9605 2900 9639
rect 2934 9636 2946 9639
rect 3694 9636 3700 9648
rect 2934 9608 3700 9636
rect 2934 9605 2946 9608
rect 2888 9599 2946 9605
rect 3694 9596 3700 9608
rect 3752 9636 3758 9648
rect 3752 9608 6914 9636
rect 3752 9596 3758 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2314 9568 2320 9580
rect 1719 9540 2320 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2464 9540 2697 9568
rect 2464 9528 2470 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3234 9568 3240 9580
rect 3099 9540 3240 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3234 9528 3240 9540
rect 3292 9568 3298 9580
rect 4614 9568 4620 9580
rect 3292 9540 4620 9568
rect 3292 9528 3298 9540
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 6886 9568 6914 9608
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 6886 9540 9229 9568
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 9217 9531 9275 9537
rect 9766 9528 9772 9580
rect 9824 9568 9830 9580
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 9824 9540 9873 9568
rect 9824 9528 9830 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 2556 9404 2789 9432
rect 2556 9392 2562 9404
rect 2777 9401 2789 9404
rect 2823 9401 2835 9435
rect 10042 9432 10048 9444
rect 10003 9404 10048 9432
rect 2777 9395 2835 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 9401 9367 9459 9373
rect 9401 9333 9413 9367
rect 9447 9364 9459 9367
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 9447 9336 11253 9364
rect 9447 9333 9459 9336
rect 9401 9327 9459 9333
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5845 9274
rect 5897 9222 5909 9274
rect 5961 9222 5973 9274
rect 6025 9222 6037 9274
rect 6089 9222 6101 9274
rect 6153 9222 9109 9274
rect 9161 9222 9173 9274
rect 9225 9222 9237 9274
rect 9289 9222 9301 9274
rect 9353 9222 9365 9274
rect 9417 9222 10856 9274
rect 1104 9200 10856 9222
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9129 2467 9163
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 2409 9123 2467 9129
rect 2424 9092 2452 9123
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 9401 9163 9459 9169
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 9447 9132 11161 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 6546 9092 6552 9104
rect 2424 9064 6552 9092
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 2464 8996 6914 9024
rect 2464 8984 2470 8996
rect 1854 8956 1860 8968
rect 1815 8928 1860 8956
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2866 8956 2872 8968
rect 2639 8928 2872 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3050 8956 3056 8968
rect 3011 8928 3056 8956
rect 3050 8916 3056 8928
rect 3108 8916 3114 8968
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 3510 8956 3516 8968
rect 3200 8928 3516 8956
rect 3200 8916 3206 8928
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 6886 8956 6914 8996
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 6886 8928 9229 8956
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9858 8956 9864 8968
rect 9819 8928 9864 8956
rect 9217 8919 9275 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 1578 8848 1584 8900
rect 1636 8888 1642 8900
rect 6454 8888 6460 8900
rect 1636 8860 6460 8888
rect 1636 8848 1642 8860
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 6178 8820 6184 8832
rect 1719 8792 6184 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 1104 8730 10856 8752
rect 1104 8678 4213 8730
rect 4265 8678 4277 8730
rect 4329 8678 4341 8730
rect 4393 8678 4405 8730
rect 4457 8678 4469 8730
rect 4521 8678 7477 8730
rect 7529 8678 7541 8730
rect 7593 8678 7605 8730
rect 7657 8678 7669 8730
rect 7721 8678 7733 8730
rect 7785 8678 10856 8730
rect 1104 8656 10856 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 2317 8619 2375 8625
rect 2317 8585 2329 8619
rect 2363 8585 2375 8619
rect 3694 8616 3700 8628
rect 3655 8588 3700 8616
rect 2317 8579 2375 8585
rect 2332 8548 2360 8579
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 6730 8548 6736 8560
rect 2332 8520 6736 8548
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8480 1455 8483
rect 1486 8480 1492 8492
rect 1443 8452 1492 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 2130 8480 2136 8492
rect 1636 8452 2136 8480
rect 1636 8440 1642 8452
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 2866 8480 2872 8492
rect 2779 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 6886 8452 9873 8480
rect 2884 8412 2912 8440
rect 3694 8412 3700 8424
rect 2884 8384 3700 8412
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 6886 8344 6914 8452
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 3099 8316 6914 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 10042 8276 10048 8288
rect 10003 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5845 8186
rect 5897 8134 5909 8186
rect 5961 8134 5973 8186
rect 6025 8134 6037 8186
rect 6089 8134 6101 8186
rect 6153 8134 9109 8186
rect 9161 8134 9173 8186
rect 9225 8134 9237 8186
rect 9289 8134 9301 8186
rect 9353 8134 9365 8186
rect 9417 8134 10856 8186
rect 1104 8112 10856 8134
rect 3970 8072 3976 8084
rect 3931 8044 3976 8072
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 3786 8004 3792 8016
rect 2832 7976 3792 8004
rect 2832 7964 2838 7976
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 2406 7936 2412 7948
rect 1719 7908 2412 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 3418 7936 3424 7948
rect 3200 7908 3424 7936
rect 3200 7896 3206 7908
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2498 7868 2504 7880
rect 1912 7840 2504 7868
rect 1912 7828 1918 7840
rect 2498 7828 2504 7840
rect 2556 7868 2562 7880
rect 2685 7871 2743 7877
rect 2685 7868 2697 7871
rect 2556 7840 2697 7868
rect 2556 7828 2562 7840
rect 2685 7837 2697 7840
rect 2731 7837 2743 7871
rect 3786 7868 3792 7880
rect 3747 7840 3792 7868
rect 2685 7831 2743 7837
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 9858 7800 9864 7812
rect 2884 7772 9864 7800
rect 2884 7741 2912 7772
rect 9858 7760 9864 7772
rect 9916 7760 9922 7812
rect 2869 7735 2927 7741
rect 2869 7701 2881 7735
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 1104 7642 10856 7664
rect 1104 7590 4213 7642
rect 4265 7590 4277 7642
rect 4329 7590 4341 7642
rect 4393 7590 4405 7642
rect 4457 7590 4469 7642
rect 4521 7590 7477 7642
rect 7529 7590 7541 7642
rect 7593 7590 7605 7642
rect 7657 7590 7669 7642
rect 7721 7590 7733 7642
rect 7785 7590 10856 7642
rect 1104 7568 10856 7590
rect 2774 7528 2780 7540
rect 2735 7500 2780 7528
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 1210 7420 1216 7472
rect 1268 7460 1274 7472
rect 1857 7463 1915 7469
rect 1857 7460 1869 7463
rect 1268 7432 1869 7460
rect 1268 7420 1274 7432
rect 1857 7429 1869 7432
rect 1903 7460 1915 7463
rect 1903 7432 3372 7460
rect 1903 7429 1915 7432
rect 1857 7423 1915 7429
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 1964 7324 1992 7355
rect 2038 7352 2044 7404
rect 2096 7392 2102 7404
rect 3344 7401 3372 7432
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2096 7364 2605 7392
rect 2096 7352 2102 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3602 7392 3608 7404
rect 3559 7364 3608 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 9858 7392 9864 7404
rect 9819 7364 9864 7392
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 3694 7324 3700 7336
rect 1964 7296 3700 7324
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 9858 7188 9864 7200
rect 3559 7160 9864 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 9858 7148 9864 7160
rect 9916 7148 9922 7200
rect 10042 7188 10048 7200
rect 10003 7160 10048 7188
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5845 7098
rect 5897 7046 5909 7098
rect 5961 7046 5973 7098
rect 6025 7046 6037 7098
rect 6089 7046 6101 7098
rect 6153 7046 9109 7098
rect 9161 7046 9173 7098
rect 9225 7046 9237 7098
rect 9289 7046 9301 7098
rect 9353 7046 9365 7098
rect 9417 7046 10856 7098
rect 1104 7024 10856 7046
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 1486 6740 1492 6792
rect 1544 6780 1550 6792
rect 2593 6783 2651 6789
rect 2593 6780 2605 6783
rect 1544 6752 2605 6780
rect 1544 6740 1550 6752
rect 2593 6749 2605 6752
rect 2639 6749 2651 6783
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 2593 6743 2651 6749
rect 6886 6752 9873 6780
rect 4062 6712 4068 6724
rect 1596 6684 4068 6712
rect 1596 6653 1624 6684
rect 4062 6672 4068 6684
rect 4120 6672 4126 6724
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 6886 6644 6914 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10042 6644 10048 6656
rect 2823 6616 6914 6644
rect 10003 6616 10048 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 1104 6554 10856 6576
rect 1104 6502 4213 6554
rect 4265 6502 4277 6554
rect 4329 6502 4341 6554
rect 4393 6502 4405 6554
rect 4457 6502 4469 6554
rect 4521 6502 7477 6554
rect 7529 6502 7541 6554
rect 7593 6502 7605 6554
rect 7657 6502 7669 6554
rect 7721 6502 7733 6554
rect 7785 6502 10856 6554
rect 1104 6480 10856 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3510 6440 3516 6452
rect 3471 6412 3516 6440
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 2958 6304 2964 6316
rect 2731 6276 2964 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3326 6304 3332 6316
rect 3287 6276 3332 6304
rect 3326 6264 3332 6276
rect 3384 6264 3390 6316
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3878 6168 3884 6180
rect 2915 6140 3884 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3878 6128 3884 6140
rect 3936 6128 3942 6180
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5845 6010
rect 5897 5958 5909 6010
rect 5961 5958 5973 6010
rect 6025 5958 6037 6010
rect 6089 5958 6101 6010
rect 6153 5958 9109 6010
rect 9161 5958 9173 6010
rect 9225 5958 9237 6010
rect 9289 5958 9301 6010
rect 9353 5958 9365 6010
rect 9417 5958 10856 6010
rect 1104 5936 10856 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1544 5868 1593 5896
rect 1544 5856 1550 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 1360 5664 1409 5692
rect 1360 5652 1366 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1578 5652 1584 5704
rect 1636 5692 1642 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 1636 5664 2329 5692
rect 1636 5652 1642 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 9861 5695 9919 5701
rect 9861 5692 9873 5695
rect 2317 5655 2375 5661
rect 6886 5664 9873 5692
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 6886 5556 6914 5664
rect 9861 5661 9873 5664
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 10042 5556 10048 5568
rect 2547 5528 6914 5556
rect 10003 5528 10048 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 1104 5466 10856 5488
rect 1104 5414 4213 5466
rect 4265 5414 4277 5466
rect 4329 5414 4341 5466
rect 4393 5414 4405 5466
rect 4457 5414 4469 5466
rect 4521 5414 7477 5466
rect 7529 5414 7541 5466
rect 7593 5414 7605 5466
rect 7657 5414 7669 5466
rect 7721 5414 7733 5466
rect 7785 5414 10856 5466
rect 1104 5392 10856 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 5534 5352 5540 5364
rect 1627 5324 5540 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 2225 5287 2283 5293
rect 2225 5253 2237 5287
rect 2271 5284 2283 5287
rect 3234 5284 3240 5296
rect 2271 5256 3240 5284
rect 2271 5253 2283 5256
rect 2225 5247 2283 5253
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1578 5216 1584 5228
rect 1443 5188 1584 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1578 5176 1584 5188
rect 1636 5176 1642 5228
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2792 5225 2820 5256
rect 3234 5244 3240 5256
rect 3292 5244 3298 5296
rect 3620 5256 4292 5284
rect 3620 5228 3648 5256
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 3418 5216 3424 5228
rect 3379 5188 3424 5216
rect 2961 5179 3019 5185
rect 2976 5148 3004 5179
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 4264 5225 4292 5256
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 9858 5216 9864 5228
rect 9819 5188 9864 5216
rect 4249 5179 4307 5185
rect 3620 5148 3648 5176
rect 2976 5120 3648 5148
rect 4080 5148 4108 5179
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 4706 5148 4712 5160
rect 4080 5120 4712 5148
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 2958 5012 2964 5024
rect 2919 4984 2964 5012
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4154 5012 4160 5024
rect 3651 4984 4160 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 7098 5012 7104 5024
rect 4295 4984 7104 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5845 4922
rect 5897 4870 5909 4922
rect 5961 4870 5973 4922
rect 6025 4870 6037 4922
rect 6089 4870 6101 4922
rect 6153 4870 9109 4922
rect 9161 4870 9173 4922
rect 9225 4870 9237 4922
rect 9289 4870 9301 4922
rect 9353 4870 9365 4922
rect 9417 4870 10856 4922
rect 1104 4848 10856 4870
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 3418 4808 3424 4820
rect 2271 4780 3424 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 9858 4808 9864 4820
rect 4212 4780 9864 4808
rect 4212 4768 4218 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4740 2835 4743
rect 4706 4740 4712 4752
rect 2823 4712 4712 4740
rect 2823 4709 2835 4712
rect 2777 4703 2835 4709
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 9766 4672 9772 4684
rect 3016 4644 9772 4672
rect 3016 4632 3022 4644
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3418 4604 3424 4616
rect 2915 4576 3424 4604
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 2240 4536 2268 4567
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 7156 4576 9873 4604
rect 7156 4564 7162 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 3786 4536 3792 4548
rect 2240 4508 3792 4536
rect 3786 4496 3792 4508
rect 3844 4496 3850 4548
rect 10042 4468 10048 4480
rect 10003 4440 10048 4468
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 1104 4378 10856 4400
rect 1104 4326 4213 4378
rect 4265 4326 4277 4378
rect 4329 4326 4341 4378
rect 4393 4326 4405 4378
rect 4457 4326 4469 4378
rect 4521 4326 7477 4378
rect 7529 4326 7541 4378
rect 7593 4326 7605 4378
rect 7657 4326 7669 4378
rect 7721 4326 7733 4378
rect 7785 4326 10856 4378
rect 1104 4304 10856 4326
rect 1946 4156 1952 4208
rect 2004 4196 2010 4208
rect 2041 4199 2099 4205
rect 2041 4196 2053 4199
rect 2004 4168 2053 4196
rect 2004 4156 2010 4168
rect 2041 4165 2053 4168
rect 2087 4165 2099 4199
rect 3602 4196 3608 4208
rect 2041 4159 2099 4165
rect 2240 4168 2452 4196
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1412 4100 1593 4128
rect 1412 3924 1440 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 2240 4060 2268 4168
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2424 4128 2452 4168
rect 3436 4168 3608 4196
rect 3436 4137 3464 4168
rect 3602 4156 3608 4168
rect 3660 4196 3666 4208
rect 3660 4168 4108 4196
rect 3660 4156 3666 4168
rect 2501 4131 2559 4137
rect 2501 4128 2513 4131
rect 2424 4100 2513 4128
rect 2317 4091 2375 4097
rect 2501 4097 2513 4100
rect 2547 4128 2559 4131
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 2547 4100 3249 4128
rect 2547 4097 2559 4100
rect 2501 4091 2559 4097
rect 3237 4097 3249 4100
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4097 3479 4131
rect 3421 4091 3479 4097
rect 1535 4032 2268 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 2332 3992 2360 4091
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 4080 4137 4108 4168
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3568 4100 3893 4128
rect 3568 4088 3574 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4097 4123 4131
rect 4065 4091 4123 4097
rect 4614 4060 4620 4072
rect 3344 4032 4620 4060
rect 3142 3992 3148 4004
rect 2332 3964 3148 3992
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3344 3924 3372 4032
rect 4614 4020 4620 4032
rect 4672 4020 4678 4072
rect 3421 3995 3479 4001
rect 3421 3961 3433 3995
rect 3467 3992 3479 3995
rect 5534 3992 5540 4004
rect 3467 3964 5540 3992
rect 3467 3961 3479 3964
rect 3421 3955 3479 3961
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 1412 3896 3372 3924
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 8018 3924 8024 3936
rect 4111 3896 8024 3924
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5845 3834
rect 5897 3782 5909 3834
rect 5961 3782 5973 3834
rect 6025 3782 6037 3834
rect 6089 3782 6101 3834
rect 6153 3782 9109 3834
rect 9161 3782 9173 3834
rect 9225 3782 9237 3834
rect 9289 3782 9301 3834
rect 9353 3782 9365 3834
rect 9417 3782 10856 3834
rect 1104 3760 10856 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 2556 3692 3801 3720
rect 2556 3680 2562 3692
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 3789 3683 3847 3689
rect 3142 3584 3148 3596
rect 2148 3556 3148 3584
rect 2148 3525 2176 3556
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2280 3488 2697 3516
rect 2280 3476 2286 3488
rect 2685 3485 2697 3488
rect 2731 3516 2743 3519
rect 3510 3516 3516 3528
rect 2731 3488 3516 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3970 3516 3976 3528
rect 3931 3488 3976 3516
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 7926 3448 7932 3460
rect 2608 3420 7932 3448
rect 2608 3389 2636 3420
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 2593 3383 2651 3389
rect 2593 3349 2605 3383
rect 2639 3349 2651 3383
rect 10042 3380 10048 3392
rect 10003 3352 10048 3380
rect 2593 3343 2651 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 1104 3290 10856 3312
rect 1104 3238 4213 3290
rect 4265 3238 4277 3290
rect 4329 3238 4341 3290
rect 4393 3238 4405 3290
rect 4457 3238 4469 3290
rect 4521 3238 7477 3290
rect 7529 3238 7541 3290
rect 7593 3238 7605 3290
rect 7657 3238 7669 3290
rect 7721 3238 7733 3290
rect 7785 3238 10856 3290
rect 1104 3216 10856 3238
rect 2222 3176 2228 3188
rect 2183 3148 2228 3176
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 3418 3176 3424 3188
rect 3379 3148 3424 3176
rect 3418 3136 3424 3148
rect 3476 3136 3482 3188
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 3752 3148 4077 3176
rect 3752 3136 3758 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 1688 3080 2452 3108
rect 1688 3049 1716 3080
rect 2424 3052 2452 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2332 2972 2360 3003
rect 2406 3000 2412 3052
rect 2464 3040 2470 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 2464 3012 2789 3040
rect 2464 3000 2470 3012
rect 2777 3009 2789 3012
rect 2823 3009 2835 3043
rect 3602 3040 3608 3052
rect 3563 3012 3608 3040
rect 2777 3003 2835 3009
rect 3602 3000 3608 3012
rect 3660 3000 3666 3052
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4212 3012 4261 3040
rect 4212 3000 4218 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 8076 3012 9137 3040
rect 8076 3000 8082 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9125 3003 9183 3009
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9824 3012 9873 3040
rect 9824 3000 9830 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 5074 2972 5080 2984
rect 2332 2944 5080 2972
rect 5074 2932 5080 2944
rect 5132 2932 5138 2984
rect 2961 2907 3019 2913
rect 2961 2873 2973 2907
rect 3007 2904 3019 2907
rect 9858 2904 9864 2916
rect 3007 2876 9864 2904
rect 3007 2873 3019 2876
rect 2961 2867 3019 2873
rect 9858 2864 9864 2876
rect 9916 2864 9922 2916
rect 1489 2839 1547 2845
rect 1489 2805 1501 2839
rect 1535 2836 1547 2839
rect 5626 2836 5632 2848
rect 1535 2808 5632 2836
rect 1535 2805 1547 2808
rect 1489 2799 1547 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 9490 2836 9496 2848
rect 9355 2808 9496 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5845 2746
rect 5897 2694 5909 2746
rect 5961 2694 5973 2746
rect 6025 2694 6037 2746
rect 6089 2694 6101 2746
rect 6153 2694 9109 2746
rect 9161 2694 9173 2746
rect 9225 2694 9237 2746
rect 9289 2694 9301 2746
rect 9353 2694 9365 2746
rect 9417 2694 10856 2746
rect 1104 2672 10856 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2372 2604 2697 2632
rect 2372 2592 2378 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 2685 2595 2743 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4433 2635 4491 2641
rect 4433 2601 4445 2635
rect 4479 2632 4491 2635
rect 4614 2632 4620 2644
rect 4479 2604 4620 2632
rect 4479 2601 4491 2604
rect 4433 2595 4491 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5074 2632 5080 2644
rect 5035 2604 5080 2632
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 2225 2567 2283 2573
rect 2225 2533 2237 2567
rect 2271 2564 2283 2567
rect 2406 2564 2412 2576
rect 2271 2536 2412 2564
rect 2271 2533 2283 2536
rect 2225 2527 2283 2533
rect 2406 2524 2412 2536
rect 2464 2524 2470 2576
rect 1394 2428 1400 2440
rect 1355 2400 1400 2428
rect 1394 2388 1400 2400
rect 1452 2388 1458 2440
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2774 2428 2780 2440
rect 2087 2400 2780 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 3970 2428 3976 2440
rect 2924 2400 2969 2428
rect 3931 2400 3976 2428
rect 2924 2388 2930 2400
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5258 2428 5264 2440
rect 5219 2400 5264 2428
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 5592 2400 9137 2428
rect 5592 2388 5598 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9858 2428 9864 2440
rect 9819 2400 9864 2428
rect 9125 2391 9183 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 1104 2202 10856 2224
rect 1104 2150 4213 2202
rect 4265 2150 4277 2202
rect 4329 2150 4341 2202
rect 4393 2150 4405 2202
rect 4457 2150 4469 2202
rect 4521 2150 7477 2202
rect 7529 2150 7541 2202
rect 7593 2150 7605 2202
rect 7657 2150 7669 2202
rect 7721 2150 7733 2202
rect 7785 2150 10856 2202
rect 1104 2128 10856 2150
rect 2866 1028 2872 1080
rect 2924 1068 2930 1080
rect 5258 1068 5264 1080
rect 2924 1040 5264 1068
rect 2924 1028 2930 1040
rect 5258 1028 5264 1040
rect 5316 1028 5322 1080
rect 2774 484 2780 536
rect 2832 524 2838 536
rect 4614 524 4620 536
rect 2832 496 4620 524
rect 2832 484 2838 496
rect 4614 484 4620 496
rect 4672 484 4678 536
<< via1 >>
rect 10968 78659 11020 78668
rect 10968 78625 10977 78659
rect 10977 78625 11011 78659
rect 11011 78625 11020 78659
rect 10968 78616 11020 78625
rect 2780 78072 2832 78124
rect 4620 78072 4672 78124
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5845 77766 5897 77818
rect 5909 77766 5961 77818
rect 5973 77766 6025 77818
rect 6037 77766 6089 77818
rect 6101 77766 6153 77818
rect 9109 77766 9161 77818
rect 9173 77766 9225 77818
rect 9237 77766 9289 77818
rect 9301 77766 9353 77818
rect 9365 77766 9417 77818
rect 1400 77571 1452 77580
rect 1400 77537 1409 77571
rect 1409 77537 1443 77571
rect 1443 77537 1452 77571
rect 1400 77528 1452 77537
rect 3608 77528 3660 77580
rect 2964 77460 3016 77512
rect 3976 77503 4028 77512
rect 3976 77469 3985 77503
rect 3985 77469 4019 77503
rect 4019 77469 4028 77503
rect 3976 77460 4028 77469
rect 4068 77460 4120 77512
rect 9404 77503 9456 77512
rect 9404 77469 9413 77503
rect 9413 77469 9447 77503
rect 9447 77469 9456 77503
rect 9404 77460 9456 77469
rect 10048 77503 10100 77512
rect 10048 77469 10057 77503
rect 10057 77469 10091 77503
rect 10091 77469 10100 77503
rect 10048 77460 10100 77469
rect 2136 77324 2188 77376
rect 3792 77367 3844 77376
rect 3792 77333 3801 77367
rect 3801 77333 3835 77367
rect 3835 77333 3844 77367
rect 3792 77324 3844 77333
rect 3884 77324 3936 77376
rect 5264 77324 5316 77376
rect 4213 77222 4265 77274
rect 4277 77222 4329 77274
rect 4341 77222 4393 77274
rect 4405 77222 4457 77274
rect 4469 77222 4521 77274
rect 7477 77222 7529 77274
rect 7541 77222 7593 77274
rect 7605 77222 7657 77274
rect 7669 77222 7721 77274
rect 7733 77222 7785 77274
rect 1400 77027 1452 77036
rect 1400 76993 1409 77027
rect 1409 76993 1443 77027
rect 1443 76993 1452 77027
rect 1400 76984 1452 76993
rect 2228 76984 2280 77036
rect 2964 76984 3016 77036
rect 3332 77027 3384 77036
rect 3332 76993 3341 77027
rect 3341 76993 3375 77027
rect 3375 76993 3384 77027
rect 3332 76984 3384 76993
rect 3424 76984 3476 77036
rect 4620 77027 4672 77036
rect 4620 76993 4629 77027
rect 4629 76993 4663 77027
rect 4663 76993 4672 77027
rect 4620 76984 4672 76993
rect 9496 76984 9548 77036
rect 5540 76848 5592 76900
rect 2412 76780 2464 76832
rect 3056 76780 3108 76832
rect 3240 76780 3292 76832
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5845 76678 5897 76730
rect 5909 76678 5961 76730
rect 5973 76678 6025 76730
rect 6037 76678 6089 76730
rect 6101 76678 6153 76730
rect 9109 76678 9161 76730
rect 9173 76678 9225 76730
rect 9237 76678 9289 76730
rect 9301 76678 9353 76730
rect 9365 76678 9417 76730
rect 112 76508 164 76560
rect 1400 76372 1452 76424
rect 1952 76372 2004 76424
rect 2228 76415 2280 76424
rect 2228 76381 2242 76415
rect 2242 76381 2276 76415
rect 2276 76381 2280 76415
rect 3148 76415 3200 76424
rect 2228 76372 2280 76381
rect 3148 76381 3157 76415
rect 3157 76381 3191 76415
rect 3191 76381 3200 76415
rect 3148 76372 3200 76381
rect 3516 76372 3568 76424
rect 10140 76415 10192 76424
rect 10140 76381 10149 76415
rect 10149 76381 10183 76415
rect 10183 76381 10192 76415
rect 10140 76372 10192 76381
rect 5264 76304 5316 76356
rect 3424 76236 3476 76288
rect 9956 76279 10008 76288
rect 9956 76245 9965 76279
rect 9965 76245 9999 76279
rect 9999 76245 10008 76279
rect 9956 76236 10008 76245
rect 4213 76134 4265 76186
rect 4277 76134 4329 76186
rect 4341 76134 4393 76186
rect 4405 76134 4457 76186
rect 4469 76134 4521 76186
rect 7477 76134 7529 76186
rect 7541 76134 7593 76186
rect 7605 76134 7657 76186
rect 7669 76134 7721 76186
rect 7733 76134 7785 76186
rect 1768 76032 1820 76084
rect 3240 76032 3292 76084
rect 3332 76032 3384 76084
rect 1492 75896 1544 75948
rect 1952 75896 2004 75948
rect 2228 75828 2280 75880
rect 3608 75939 3660 75948
rect 3608 75905 3617 75939
rect 3617 75905 3651 75939
rect 3651 75905 3660 75939
rect 3608 75896 3660 75905
rect 10232 75828 10284 75880
rect 3240 75760 3292 75812
rect 3516 75760 3568 75812
rect 3976 75692 4028 75744
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5845 75590 5897 75642
rect 5909 75590 5961 75642
rect 5973 75590 6025 75642
rect 6037 75590 6089 75642
rect 6101 75590 6153 75642
rect 9109 75590 9161 75642
rect 9173 75590 9225 75642
rect 9237 75590 9289 75642
rect 9301 75590 9353 75642
rect 9365 75590 9417 75642
rect 8300 75420 8352 75472
rect 1952 75284 2004 75336
rect 3884 75352 3936 75404
rect 2228 75327 2280 75336
rect 2228 75293 2242 75327
rect 2242 75293 2276 75327
rect 2276 75293 2280 75327
rect 3148 75327 3200 75336
rect 2228 75284 2280 75293
rect 3148 75293 3157 75327
rect 3157 75293 3191 75327
rect 3191 75293 3200 75327
rect 3148 75284 3200 75293
rect 9956 75284 10008 75336
rect 10140 75327 10192 75336
rect 10140 75293 10149 75327
rect 10149 75293 10183 75327
rect 10183 75293 10192 75327
rect 10140 75284 10192 75293
rect 2964 75191 3016 75200
rect 2964 75157 2973 75191
rect 2973 75157 3007 75191
rect 3007 75157 3016 75191
rect 2964 75148 3016 75157
rect 9956 75191 10008 75200
rect 9956 75157 9965 75191
rect 9965 75157 9999 75191
rect 9999 75157 10008 75191
rect 9956 75148 10008 75157
rect 4213 75046 4265 75098
rect 4277 75046 4329 75098
rect 4341 75046 4393 75098
rect 4405 75046 4457 75098
rect 4469 75046 4521 75098
rect 7477 75046 7529 75098
rect 7541 75046 7593 75098
rect 7605 75046 7657 75098
rect 7669 75046 7721 75098
rect 7733 75046 7785 75098
rect 3792 74876 3844 74928
rect 1400 74851 1452 74860
rect 1400 74817 1409 74851
rect 1409 74817 1443 74851
rect 1443 74817 1452 74851
rect 1400 74808 1452 74817
rect 1676 74808 1728 74860
rect 2228 74808 2280 74860
rect 3148 74808 3200 74860
rect 9956 74740 10008 74792
rect 1584 74647 1636 74656
rect 1584 74613 1593 74647
rect 1593 74613 1627 74647
rect 1627 74613 1636 74647
rect 1584 74604 1636 74613
rect 5632 74604 5684 74656
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5845 74502 5897 74554
rect 5909 74502 5961 74554
rect 5973 74502 6025 74554
rect 6037 74502 6089 74554
rect 6101 74502 6153 74554
rect 9109 74502 9161 74554
rect 9173 74502 9225 74554
rect 9237 74502 9289 74554
rect 9301 74502 9353 74554
rect 9365 74502 9417 74554
rect 1400 74239 1452 74248
rect 1400 74205 1409 74239
rect 1409 74205 1443 74239
rect 1443 74205 1452 74239
rect 1400 74196 1452 74205
rect 10140 74239 10192 74248
rect 10140 74205 10149 74239
rect 10149 74205 10183 74239
rect 10183 74205 10192 74239
rect 10140 74196 10192 74205
rect 1492 74060 1544 74112
rect 9956 74103 10008 74112
rect 9956 74069 9965 74103
rect 9965 74069 9999 74103
rect 9999 74069 10008 74103
rect 9956 74060 10008 74069
rect 4213 73958 4265 74010
rect 4277 73958 4329 74010
rect 4341 73958 4393 74010
rect 4405 73958 4457 74010
rect 4469 73958 4521 74010
rect 7477 73958 7529 74010
rect 7541 73958 7593 74010
rect 7605 73958 7657 74010
rect 7669 73958 7721 74010
rect 7733 73958 7785 74010
rect 2964 73788 3016 73840
rect 1676 73763 1728 73772
rect 1676 73729 1680 73763
rect 1680 73729 1714 73763
rect 1714 73729 1728 73763
rect 1676 73720 1728 73729
rect 1952 73720 2004 73772
rect 2228 73720 2280 73772
rect 2780 73720 2832 73772
rect 10140 73763 10192 73772
rect 10140 73729 10149 73763
rect 10149 73729 10183 73763
rect 10183 73729 10192 73763
rect 10140 73720 10192 73729
rect 9864 73652 9916 73704
rect 572 73516 624 73568
rect 1952 73516 2004 73568
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5845 73414 5897 73466
rect 5909 73414 5961 73466
rect 5973 73414 6025 73466
rect 6037 73414 6089 73466
rect 6101 73414 6153 73466
rect 9109 73414 9161 73466
rect 9173 73414 9225 73466
rect 9237 73414 9289 73466
rect 9301 73414 9353 73466
rect 9365 73414 9417 73466
rect 1676 73151 1728 73160
rect 1676 73117 1680 73151
rect 1680 73117 1714 73151
rect 1714 73117 1728 73151
rect 1676 73108 1728 73117
rect 1860 73083 1912 73092
rect 1860 73049 1869 73083
rect 1869 73049 1903 73083
rect 1903 73049 1912 73083
rect 1860 73040 1912 73049
rect 2228 73176 2280 73228
rect 2964 73176 3016 73228
rect 3148 73176 3200 73228
rect 2780 73108 2832 73160
rect 4068 73040 4120 73092
rect 2228 72972 2280 73024
rect 2504 72972 2556 73024
rect 4213 72870 4265 72922
rect 4277 72870 4329 72922
rect 4341 72870 4393 72922
rect 4405 72870 4457 72922
rect 4469 72870 4521 72922
rect 7477 72870 7529 72922
rect 7541 72870 7593 72922
rect 7605 72870 7657 72922
rect 7669 72870 7721 72922
rect 7733 72870 7785 72922
rect 1860 72768 1912 72820
rect 3332 72768 3384 72820
rect 9956 72700 10008 72752
rect 1400 72675 1452 72684
rect 1400 72641 1409 72675
rect 1409 72641 1443 72675
rect 1443 72641 1452 72675
rect 1400 72632 1452 72641
rect 1676 72632 1728 72684
rect 2320 72632 2372 72684
rect 2964 72632 3016 72684
rect 10140 72675 10192 72684
rect 10140 72641 10149 72675
rect 10149 72641 10183 72675
rect 10183 72641 10192 72675
rect 10140 72632 10192 72641
rect 3056 72564 3108 72616
rect 4068 72564 4120 72616
rect 9956 72564 10008 72616
rect 2228 72496 2280 72548
rect 8392 72496 8444 72548
rect 1676 72428 1728 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5845 72326 5897 72378
rect 5909 72326 5961 72378
rect 5973 72326 6025 72378
rect 6037 72326 6089 72378
rect 6101 72326 6153 72378
rect 9109 72326 9161 72378
rect 9173 72326 9225 72378
rect 9237 72326 9289 72378
rect 9301 72326 9353 72378
rect 9365 72326 9417 72378
rect 9956 72267 10008 72276
rect 9956 72233 9965 72267
rect 9965 72233 9999 72267
rect 9999 72233 10008 72267
rect 9956 72224 10008 72233
rect 1216 72020 1268 72072
rect 2044 72063 2096 72072
rect 2044 72029 2053 72063
rect 2053 72029 2087 72063
rect 2087 72029 2096 72063
rect 2044 72020 2096 72029
rect 10140 72063 10192 72072
rect 10140 72029 10149 72063
rect 10149 72029 10183 72063
rect 10183 72029 10192 72063
rect 10140 72020 10192 72029
rect 1492 71884 1544 71936
rect 2320 71884 2372 71936
rect 4213 71782 4265 71834
rect 4277 71782 4329 71834
rect 4341 71782 4393 71834
rect 4405 71782 4457 71834
rect 4469 71782 4521 71834
rect 7477 71782 7529 71834
rect 7541 71782 7593 71834
rect 7605 71782 7657 71834
rect 7669 71782 7721 71834
rect 7733 71782 7785 71834
rect 2044 71680 2096 71732
rect 2228 71680 2280 71732
rect 9864 71680 9916 71732
rect 1308 71544 1360 71596
rect 2228 71587 2280 71596
rect 2228 71553 2237 71587
rect 2237 71553 2271 71587
rect 2271 71553 2280 71587
rect 2228 71544 2280 71553
rect 10140 71587 10192 71596
rect 10140 71553 10149 71587
rect 10149 71553 10183 71587
rect 10183 71553 10192 71587
rect 10140 71544 10192 71553
rect 1860 71340 1912 71392
rect 2228 71340 2280 71392
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5845 71238 5897 71290
rect 5909 71238 5961 71290
rect 5973 71238 6025 71290
rect 6037 71238 6089 71290
rect 6101 71238 6153 71290
rect 9109 71238 9161 71290
rect 9173 71238 9225 71290
rect 9237 71238 9289 71290
rect 9301 71238 9353 71290
rect 9365 71238 9417 71290
rect 5080 71068 5132 71120
rect 2044 71000 2096 71052
rect 1400 70975 1452 70984
rect 1400 70941 1409 70975
rect 1409 70941 1443 70975
rect 1443 70941 1452 70975
rect 1400 70932 1452 70941
rect 2412 70975 2464 70984
rect 1216 70864 1268 70916
rect 2412 70941 2421 70975
rect 2421 70941 2455 70975
rect 2455 70941 2464 70975
rect 2412 70932 2464 70941
rect 2596 70975 2648 70984
rect 2596 70941 2610 70975
rect 2610 70941 2644 70975
rect 2644 70941 2648 70975
rect 2596 70932 2648 70941
rect 2044 70796 2096 70848
rect 2964 70796 3016 70848
rect 4213 70694 4265 70746
rect 4277 70694 4329 70746
rect 4341 70694 4393 70746
rect 4405 70694 4457 70746
rect 4469 70694 4521 70746
rect 7477 70694 7529 70746
rect 7541 70694 7593 70746
rect 7605 70694 7657 70746
rect 7669 70694 7721 70746
rect 7733 70694 7785 70746
rect 1768 70592 1820 70644
rect 2412 70592 2464 70644
rect 1308 70456 1360 70508
rect 1768 70499 1820 70508
rect 1768 70465 1782 70499
rect 1782 70465 1816 70499
rect 1816 70465 1820 70499
rect 1768 70456 1820 70465
rect 2596 70456 2648 70508
rect 2964 70456 3016 70508
rect 5724 70388 5776 70440
rect 10140 70320 10192 70372
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5845 70150 5897 70202
rect 5909 70150 5961 70202
rect 5973 70150 6025 70202
rect 6037 70150 6089 70202
rect 6101 70150 6153 70202
rect 9109 70150 9161 70202
rect 9173 70150 9225 70202
rect 9237 70150 9289 70202
rect 9301 70150 9353 70202
rect 9365 70150 9417 70202
rect 3608 69980 3660 70032
rect 1400 69887 1452 69896
rect 1400 69853 1409 69887
rect 1409 69853 1443 69887
rect 1443 69853 1452 69887
rect 1400 69844 1452 69853
rect 1584 69887 1636 69896
rect 1584 69853 1593 69887
rect 1593 69853 1627 69887
rect 1627 69853 1636 69887
rect 1584 69844 1636 69853
rect 1768 69887 1820 69896
rect 1768 69853 1782 69887
rect 1782 69853 1816 69887
rect 1816 69853 1820 69887
rect 1768 69844 1820 69853
rect 3056 69844 3108 69896
rect 10140 69887 10192 69896
rect 10140 69853 10149 69887
rect 10149 69853 10183 69887
rect 10183 69853 10192 69887
rect 10140 69844 10192 69853
rect 1584 69708 1636 69760
rect 2228 69708 2280 69760
rect 2596 69708 2648 69760
rect 4213 69606 4265 69658
rect 4277 69606 4329 69658
rect 4341 69606 4393 69658
rect 4405 69606 4457 69658
rect 4469 69606 4521 69658
rect 7477 69606 7529 69658
rect 7541 69606 7593 69658
rect 7605 69606 7657 69658
rect 7669 69606 7721 69658
rect 7733 69606 7785 69658
rect 1400 69504 1452 69556
rect 1952 69436 2004 69488
rect 1308 69300 1360 69352
rect 1768 69411 1820 69420
rect 1768 69377 1782 69411
rect 1782 69377 1816 69411
rect 1816 69377 1820 69411
rect 1768 69368 1820 69377
rect 2964 69368 3016 69420
rect 3332 69411 3384 69420
rect 3332 69377 3341 69411
rect 3341 69377 3375 69411
rect 3375 69377 3384 69411
rect 3332 69368 3384 69377
rect 9956 69300 10008 69352
rect 2596 69232 2648 69284
rect 1216 69164 1268 69216
rect 2136 69164 2188 69216
rect 3516 69164 3568 69216
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5845 69062 5897 69114
rect 5909 69062 5961 69114
rect 5973 69062 6025 69114
rect 6037 69062 6089 69114
rect 6101 69062 6153 69114
rect 9109 69062 9161 69114
rect 9173 69062 9225 69114
rect 9237 69062 9289 69114
rect 9301 69062 9353 69114
rect 9365 69062 9417 69114
rect 1400 68960 1452 69012
rect 1952 68960 2004 69012
rect 9956 69003 10008 69012
rect 9956 68969 9965 69003
rect 9965 68969 9999 69003
rect 9999 68969 10008 69003
rect 9956 68960 10008 68969
rect 2596 68892 2648 68944
rect 1768 68824 1820 68876
rect 1400 68799 1452 68808
rect 1400 68765 1409 68799
rect 1409 68765 1443 68799
rect 1443 68765 1452 68799
rect 1400 68756 1452 68765
rect 2872 68799 2924 68808
rect 2872 68765 2881 68799
rect 2881 68765 2915 68799
rect 2915 68765 2924 68799
rect 2872 68756 2924 68765
rect 10140 68799 10192 68808
rect 10140 68765 10149 68799
rect 10149 68765 10183 68799
rect 10183 68765 10192 68799
rect 10140 68756 10192 68765
rect 3424 68688 3476 68740
rect 1768 68620 1820 68672
rect 7012 68620 7064 68672
rect 4213 68518 4265 68570
rect 4277 68518 4329 68570
rect 4341 68518 4393 68570
rect 4405 68518 4457 68570
rect 4469 68518 4521 68570
rect 7477 68518 7529 68570
rect 7541 68518 7593 68570
rect 7605 68518 7657 68570
rect 7669 68518 7721 68570
rect 7733 68518 7785 68570
rect 1584 68416 1636 68468
rect 1032 68280 1084 68332
rect 1308 68212 1360 68264
rect 1676 68144 1728 68196
rect 1952 68348 2004 68400
rect 2780 68280 2832 68332
rect 3056 68323 3108 68332
rect 3056 68289 3070 68323
rect 3070 68289 3104 68323
rect 3104 68289 3108 68323
rect 10140 68323 10192 68332
rect 3056 68280 3108 68289
rect 10140 68289 10149 68323
rect 10149 68289 10183 68323
rect 10183 68289 10192 68323
rect 10140 68280 10192 68289
rect 2596 68212 2648 68264
rect 5172 68076 5224 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5845 67974 5897 68026
rect 5909 67974 5961 68026
rect 5973 67974 6025 68026
rect 6037 67974 6089 68026
rect 6101 67974 6153 68026
rect 9109 67974 9161 68026
rect 9173 67974 9225 68026
rect 9237 67974 9289 68026
rect 9301 67974 9353 68026
rect 9365 67974 9417 68026
rect 1124 67736 1176 67788
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 4213 67430 4265 67482
rect 4277 67430 4329 67482
rect 4341 67430 4393 67482
rect 4405 67430 4457 67482
rect 4469 67430 4521 67482
rect 7477 67430 7529 67482
rect 7541 67430 7593 67482
rect 7605 67430 7657 67482
rect 7669 67430 7721 67482
rect 7733 67430 7785 67482
rect 388 67192 440 67244
rect 10140 67235 10192 67244
rect 10140 67201 10149 67235
rect 10149 67201 10183 67235
rect 10183 67201 10192 67235
rect 10140 67192 10192 67201
rect 1400 67167 1452 67176
rect 1400 67133 1409 67167
rect 1409 67133 1443 67167
rect 1443 67133 1452 67167
rect 1400 67124 1452 67133
rect 9956 67031 10008 67040
rect 9956 66997 9965 67031
rect 9965 66997 9999 67031
rect 9999 66997 10008 67031
rect 9956 66988 10008 66997
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5845 66886 5897 66938
rect 5909 66886 5961 66938
rect 5973 66886 6025 66938
rect 6037 66886 6089 66938
rect 6101 66886 6153 66938
rect 9109 66886 9161 66938
rect 9173 66886 9225 66938
rect 9237 66886 9289 66938
rect 9301 66886 9353 66938
rect 9365 66886 9417 66938
rect 3240 66716 3292 66768
rect 3792 66716 3844 66768
rect 1400 66623 1452 66632
rect 1400 66589 1409 66623
rect 1409 66589 1443 66623
rect 1443 66589 1452 66623
rect 1400 66580 1452 66589
rect 1860 66580 1912 66632
rect 3240 66580 3292 66632
rect 10140 66623 10192 66632
rect 10140 66589 10149 66623
rect 10149 66589 10183 66623
rect 10183 66589 10192 66623
rect 10140 66580 10192 66589
rect 2320 66512 2372 66564
rect 3148 66512 3200 66564
rect 2228 66444 2280 66496
rect 2964 66444 3016 66496
rect 9864 66444 9916 66496
rect 4213 66342 4265 66394
rect 4277 66342 4329 66394
rect 4341 66342 4393 66394
rect 4405 66342 4457 66394
rect 4469 66342 4521 66394
rect 7477 66342 7529 66394
rect 7541 66342 7593 66394
rect 7605 66342 7657 66394
rect 7669 66342 7721 66394
rect 7733 66342 7785 66394
rect 1308 66240 1360 66292
rect 1676 66240 1728 66292
rect 1584 66215 1636 66224
rect 1584 66181 1593 66215
rect 1593 66181 1627 66215
rect 1627 66181 1636 66215
rect 1584 66172 1636 66181
rect 1676 66147 1728 66156
rect 1676 66113 1685 66147
rect 1685 66113 1719 66147
rect 1719 66113 1728 66147
rect 1676 66104 1728 66113
rect 2228 66036 2280 66088
rect 2872 66240 2924 66292
rect 2596 66172 2648 66224
rect 9956 66172 10008 66224
rect 2504 66147 2556 66156
rect 2504 66113 2513 66147
rect 2513 66113 2547 66147
rect 2547 66113 2556 66147
rect 2504 66104 2556 66113
rect 3056 66104 3108 66156
rect 10140 66147 10192 66156
rect 10140 66113 10149 66147
rect 10149 66113 10183 66147
rect 10183 66113 10192 66147
rect 10140 66104 10192 66113
rect 7104 65968 7156 66020
rect 7196 65968 7248 66020
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5845 65798 5897 65850
rect 5909 65798 5961 65850
rect 5973 65798 6025 65850
rect 6037 65798 6089 65850
rect 6101 65798 6153 65850
rect 9109 65798 9161 65850
rect 9173 65798 9225 65850
rect 9237 65798 9289 65850
rect 9301 65798 9353 65850
rect 9365 65798 9417 65850
rect 1768 65628 1820 65680
rect 1676 65560 1728 65612
rect 1952 65560 2004 65612
rect 1400 65535 1452 65544
rect 1400 65501 1409 65535
rect 1409 65501 1443 65535
rect 1443 65501 1452 65535
rect 1400 65492 1452 65501
rect 3148 65628 3200 65680
rect 7104 65696 7156 65748
rect 5908 65628 5960 65680
rect 9864 65560 9916 65612
rect 2688 65535 2740 65544
rect 2688 65501 2697 65535
rect 2697 65501 2731 65535
rect 2731 65501 2740 65535
rect 2688 65492 2740 65501
rect 3056 65424 3108 65476
rect 3148 65424 3200 65476
rect 1768 65356 1820 65408
rect 3332 65356 3384 65408
rect 4213 65254 4265 65306
rect 4277 65254 4329 65306
rect 4341 65254 4393 65306
rect 4405 65254 4457 65306
rect 4469 65254 4521 65306
rect 7477 65254 7529 65306
rect 7541 65254 7593 65306
rect 7605 65254 7657 65306
rect 7669 65254 7721 65306
rect 7733 65254 7785 65306
rect 6828 65152 6880 65204
rect 2044 65016 2096 65068
rect 2228 65016 2280 65068
rect 3056 65016 3108 65068
rect 3424 65016 3476 65068
rect 10140 65059 10192 65068
rect 10140 65025 10149 65059
rect 10149 65025 10183 65059
rect 10183 65025 10192 65059
rect 10140 65016 10192 65025
rect 3884 64923 3936 64932
rect 3884 64889 3893 64923
rect 3893 64889 3927 64923
rect 3927 64889 3936 64923
rect 3884 64880 3936 64889
rect 2136 64812 2188 64864
rect 3424 64812 3476 64864
rect 3608 64812 3660 64864
rect 6368 64812 6420 64864
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5845 64710 5897 64762
rect 5909 64710 5961 64762
rect 5973 64710 6025 64762
rect 6037 64710 6089 64762
rect 6101 64710 6153 64762
rect 9109 64710 9161 64762
rect 9173 64710 9225 64762
rect 9237 64710 9289 64762
rect 9301 64710 9353 64762
rect 9365 64710 9417 64762
rect 6920 64540 6972 64592
rect 1492 64404 1544 64456
rect 2044 64404 2096 64456
rect 2228 64404 2280 64456
rect 10140 64447 10192 64456
rect 10140 64413 10149 64447
rect 10149 64413 10183 64447
rect 10183 64413 10192 64447
rect 10140 64404 10192 64413
rect 6368 64336 6420 64388
rect 2780 64268 2832 64320
rect 9956 64311 10008 64320
rect 9956 64277 9965 64311
rect 9965 64277 9999 64311
rect 9999 64277 10008 64311
rect 9956 64268 10008 64277
rect 4213 64166 4265 64218
rect 4277 64166 4329 64218
rect 4341 64166 4393 64218
rect 4405 64166 4457 64218
rect 4469 64166 4521 64218
rect 7477 64166 7529 64218
rect 7541 64166 7593 64218
rect 7605 64166 7657 64218
rect 7669 64166 7721 64218
rect 7733 64166 7785 64218
rect 2228 63996 2280 64048
rect 3700 63928 3752 63980
rect 4620 63860 4672 63912
rect 1400 63724 1452 63776
rect 2228 63767 2280 63776
rect 2228 63733 2237 63767
rect 2237 63733 2271 63767
rect 2271 63733 2280 63767
rect 2228 63724 2280 63733
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5845 63622 5897 63674
rect 5909 63622 5961 63674
rect 5973 63622 6025 63674
rect 6037 63622 6089 63674
rect 6101 63622 6153 63674
rect 9109 63622 9161 63674
rect 9173 63622 9225 63674
rect 9237 63622 9289 63674
rect 9301 63622 9353 63674
rect 9365 63622 9417 63674
rect 2872 63452 2924 63504
rect 940 63316 992 63368
rect 2044 63316 2096 63368
rect 2504 63316 2556 63368
rect 10140 63359 10192 63368
rect 10140 63325 10149 63359
rect 10149 63325 10183 63359
rect 10183 63325 10192 63359
rect 10140 63316 10192 63325
rect 1492 63223 1544 63232
rect 1492 63189 1501 63223
rect 1501 63189 1535 63223
rect 1535 63189 1544 63223
rect 1492 63180 1544 63189
rect 3056 63223 3108 63232
rect 3056 63189 3065 63223
rect 3065 63189 3099 63223
rect 3099 63189 3108 63223
rect 3056 63180 3108 63189
rect 9864 63180 9916 63232
rect 4213 63078 4265 63130
rect 4277 63078 4329 63130
rect 4341 63078 4393 63130
rect 4405 63078 4457 63130
rect 4469 63078 4521 63130
rect 7477 63078 7529 63130
rect 7541 63078 7593 63130
rect 7605 63078 7657 63130
rect 7669 63078 7721 63130
rect 7733 63078 7785 63130
rect 1584 62951 1636 62960
rect 1584 62917 1593 62951
rect 1593 62917 1627 62951
rect 1627 62917 1636 62951
rect 1584 62908 1636 62917
rect 9956 62908 10008 62960
rect 2136 62840 2188 62892
rect 3332 62840 3384 62892
rect 10140 62883 10192 62892
rect 10140 62849 10149 62883
rect 10149 62849 10183 62883
rect 10183 62849 10192 62883
rect 10140 62840 10192 62849
rect 8484 62704 8536 62756
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5845 62534 5897 62586
rect 5909 62534 5961 62586
rect 5973 62534 6025 62586
rect 6037 62534 6089 62586
rect 6101 62534 6153 62586
rect 9109 62534 9161 62586
rect 9173 62534 9225 62586
rect 9237 62534 9289 62586
rect 9301 62534 9353 62586
rect 9365 62534 9417 62586
rect 1400 62296 1452 62348
rect 2044 62296 2096 62348
rect 2412 62296 2464 62348
rect 848 62228 900 62280
rect 2964 62271 3016 62280
rect 2964 62237 2973 62271
rect 2973 62237 3007 62271
rect 3007 62237 3016 62271
rect 2964 62228 3016 62237
rect 10140 62271 10192 62280
rect 10140 62237 10149 62271
rect 10149 62237 10183 62271
rect 10183 62237 10192 62271
rect 10140 62228 10192 62237
rect 1400 62092 1452 62144
rect 9772 62092 9824 62144
rect 4213 61990 4265 62042
rect 4277 61990 4329 62042
rect 4341 61990 4393 62042
rect 4405 61990 4457 62042
rect 4469 61990 4521 62042
rect 7477 61990 7529 62042
rect 7541 61990 7593 62042
rect 7605 61990 7657 62042
rect 7669 61990 7721 62042
rect 7733 61990 7785 62042
rect 204 61752 256 61804
rect 2044 61752 2096 61804
rect 1492 61684 1544 61736
rect 1492 61591 1544 61600
rect 1492 61557 1501 61591
rect 1501 61557 1535 61591
rect 1535 61557 1544 61591
rect 1492 61548 1544 61557
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5845 61446 5897 61498
rect 5909 61446 5961 61498
rect 5973 61446 6025 61498
rect 6037 61446 6089 61498
rect 6101 61446 6153 61498
rect 9109 61446 9161 61498
rect 9173 61446 9225 61498
rect 9237 61446 9289 61498
rect 9301 61446 9353 61498
rect 9365 61446 9417 61498
rect 4068 61344 4120 61396
rect 2964 61276 3016 61328
rect 3608 61276 3660 61328
rect 3792 61208 3844 61260
rect 3332 61140 3384 61192
rect 3884 61140 3936 61192
rect 10140 61183 10192 61192
rect 10140 61149 10149 61183
rect 10149 61149 10183 61183
rect 10183 61149 10192 61183
rect 10140 61140 10192 61149
rect 1400 61004 1452 61056
rect 3148 61004 3200 61056
rect 9956 61047 10008 61056
rect 9956 61013 9965 61047
rect 9965 61013 9999 61047
rect 9999 61013 10008 61047
rect 9956 61004 10008 61013
rect 4213 60902 4265 60954
rect 4277 60902 4329 60954
rect 4341 60902 4393 60954
rect 4405 60902 4457 60954
rect 4469 60902 4521 60954
rect 7477 60902 7529 60954
rect 7541 60902 7593 60954
rect 7605 60902 7657 60954
rect 7669 60902 7721 60954
rect 7733 60902 7785 60954
rect 1676 60775 1728 60784
rect 1676 60741 1685 60775
rect 1685 60741 1719 60775
rect 1719 60741 1728 60775
rect 1676 60732 1728 60741
rect 2136 60800 2188 60852
rect 2596 60800 2648 60852
rect 1676 60596 1728 60648
rect 2228 60596 2280 60648
rect 9864 60732 9916 60784
rect 10140 60707 10192 60716
rect 10140 60673 10149 60707
rect 10149 60673 10183 60707
rect 10183 60673 10192 60707
rect 10140 60664 10192 60673
rect 2780 60571 2832 60580
rect 2780 60537 2789 60571
rect 2789 60537 2823 60571
rect 2823 60537 2832 60571
rect 2780 60528 2832 60537
rect 480 60460 532 60512
rect 1216 60460 1268 60512
rect 6368 60460 6420 60512
rect 9956 60503 10008 60512
rect 9956 60469 9965 60503
rect 9965 60469 9999 60503
rect 9999 60469 10008 60503
rect 9956 60460 10008 60469
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5845 60358 5897 60410
rect 5909 60358 5961 60410
rect 5973 60358 6025 60410
rect 6037 60358 6089 60410
rect 6101 60358 6153 60410
rect 9109 60358 9161 60410
rect 9173 60358 9225 60410
rect 9237 60358 9289 60410
rect 9301 60358 9353 60410
rect 9365 60358 9417 60410
rect 2504 60256 2556 60308
rect 1216 60188 1268 60240
rect 1676 60052 1728 60104
rect 2596 60052 2648 60104
rect 9864 59984 9916 60036
rect 3516 59916 3568 59968
rect 4213 59814 4265 59866
rect 4277 59814 4329 59866
rect 4341 59814 4393 59866
rect 4405 59814 4457 59866
rect 4469 59814 4521 59866
rect 7477 59814 7529 59866
rect 7541 59814 7593 59866
rect 7605 59814 7657 59866
rect 7669 59814 7721 59866
rect 7733 59814 7785 59866
rect 1676 59712 1728 59764
rect 2320 59687 2372 59696
rect 2320 59653 2329 59687
rect 2329 59653 2363 59687
rect 2363 59653 2372 59687
rect 2320 59644 2372 59653
rect 9772 59644 9824 59696
rect 2596 59619 2648 59628
rect 2596 59585 2599 59619
rect 2599 59585 2648 59619
rect 2596 59576 2648 59585
rect 2688 59576 2740 59628
rect 10140 59619 10192 59628
rect 10140 59585 10149 59619
rect 10149 59585 10183 59619
rect 10183 59585 10192 59619
rect 10140 59576 10192 59585
rect 2320 59508 2372 59560
rect 4988 59508 5040 59560
rect 3056 59440 3108 59492
rect 1492 59415 1544 59424
rect 1492 59381 1501 59415
rect 1501 59381 1535 59415
rect 1535 59381 1544 59415
rect 1492 59372 1544 59381
rect 3240 59372 3292 59424
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5845 59270 5897 59322
rect 5909 59270 5961 59322
rect 5973 59270 6025 59322
rect 6037 59270 6089 59322
rect 6101 59270 6153 59322
rect 9109 59270 9161 59322
rect 9173 59270 9225 59322
rect 9237 59270 9289 59322
rect 9301 59270 9353 59322
rect 9365 59270 9417 59322
rect 1400 59168 1452 59220
rect 1584 59100 1636 59152
rect 1676 59032 1728 59084
rect 1584 59007 1636 59016
rect 1308 58828 1360 58880
rect 1584 58973 1593 59007
rect 1593 58973 1627 59007
rect 1627 58973 1636 59007
rect 1584 58964 1636 58973
rect 2320 58964 2372 59016
rect 3792 58964 3844 59016
rect 9956 58964 10008 59016
rect 10140 59007 10192 59016
rect 10140 58973 10149 59007
rect 10149 58973 10183 59007
rect 10183 58973 10192 59007
rect 10140 58964 10192 58973
rect 9956 58871 10008 58880
rect 9956 58837 9965 58871
rect 9965 58837 9999 58871
rect 9999 58837 10008 58871
rect 9956 58828 10008 58837
rect 4213 58726 4265 58778
rect 4277 58726 4329 58778
rect 4341 58726 4393 58778
rect 4405 58726 4457 58778
rect 4469 58726 4521 58778
rect 7477 58726 7529 58778
rect 7541 58726 7593 58778
rect 7605 58726 7657 58778
rect 7669 58726 7721 58778
rect 7733 58726 7785 58778
rect 664 58624 716 58676
rect 1676 58531 1728 58540
rect 1676 58497 1725 58531
rect 1725 58497 1728 58531
rect 1952 58531 2004 58540
rect 1676 58488 1728 58497
rect 1952 58497 1961 58531
rect 1961 58497 1995 58531
rect 1995 58497 2004 58531
rect 1952 58488 2004 58497
rect 1308 58420 1360 58472
rect 10140 58463 10192 58472
rect 10140 58429 10149 58463
rect 10149 58429 10183 58463
rect 10183 58429 10192 58463
rect 10140 58420 10192 58429
rect 8576 58352 8628 58404
rect 2412 58284 2464 58336
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5845 58182 5897 58234
rect 5909 58182 5961 58234
rect 5973 58182 6025 58234
rect 6037 58182 6089 58234
rect 6101 58182 6153 58234
rect 9109 58182 9161 58234
rect 9173 58182 9225 58234
rect 9237 58182 9289 58234
rect 9301 58182 9353 58234
rect 9365 58182 9417 58234
rect 1308 57944 1360 57996
rect 2412 58012 2464 58064
rect 3516 58012 3568 58064
rect 4068 58012 4120 58064
rect 1676 57944 1728 57996
rect 1952 57919 2004 57928
rect 1952 57885 1955 57919
rect 1955 57885 2004 57919
rect 1952 57876 2004 57885
rect 2596 57919 2648 57928
rect 2596 57885 2605 57919
rect 2605 57885 2639 57919
rect 2639 57885 2648 57919
rect 2596 57876 2648 57885
rect 3056 57876 3108 57928
rect 3884 57919 3936 57928
rect 3884 57885 3893 57919
rect 3893 57885 3927 57919
rect 3927 57885 3936 57919
rect 3884 57876 3936 57885
rect 4068 57876 4120 57928
rect 9956 57808 10008 57860
rect 2320 57740 2372 57792
rect 2780 57783 2832 57792
rect 2780 57749 2789 57783
rect 2789 57749 2823 57783
rect 2823 57749 2832 57783
rect 2780 57740 2832 57749
rect 3240 57740 3292 57792
rect 3884 57740 3936 57792
rect 4213 57638 4265 57690
rect 4277 57638 4329 57690
rect 4341 57638 4393 57690
rect 4405 57638 4457 57690
rect 4469 57638 4521 57690
rect 7477 57638 7529 57690
rect 7541 57638 7593 57690
rect 7605 57638 7657 57690
rect 7669 57638 7721 57690
rect 7733 57638 7785 57690
rect 112 57536 164 57588
rect 2596 57536 2648 57588
rect 3332 57536 3384 57588
rect 4896 57468 4948 57520
rect 1492 57239 1544 57248
rect 1492 57205 1501 57239
rect 1501 57205 1535 57239
rect 1535 57205 1544 57239
rect 1492 57196 1544 57205
rect 3240 57400 3292 57452
rect 3332 57332 3384 57384
rect 10140 57375 10192 57384
rect 10140 57341 10149 57375
rect 10149 57341 10183 57375
rect 10183 57341 10192 57375
rect 10140 57332 10192 57341
rect 2228 57307 2280 57316
rect 2228 57273 2237 57307
rect 2237 57273 2271 57307
rect 2271 57273 2280 57307
rect 2228 57264 2280 57273
rect 5356 57196 5408 57248
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5845 57094 5897 57146
rect 5909 57094 5961 57146
rect 5973 57094 6025 57146
rect 6037 57094 6089 57146
rect 6101 57094 6153 57146
rect 9109 57094 9161 57146
rect 9173 57094 9225 57146
rect 9237 57094 9289 57146
rect 9301 57094 9353 57146
rect 9365 57094 9417 57146
rect 2964 56992 3016 57044
rect 2412 56924 2464 56976
rect 2596 56924 2648 56976
rect 756 56788 808 56840
rect 2412 56831 2464 56840
rect 2412 56797 2421 56831
rect 2421 56797 2455 56831
rect 2455 56797 2464 56831
rect 2412 56788 2464 56797
rect 3332 56788 3384 56840
rect 6644 56856 6696 56908
rect 3516 56720 3568 56772
rect 4068 56788 4120 56840
rect 10140 56831 10192 56840
rect 10140 56797 10149 56831
rect 10149 56797 10183 56831
rect 10183 56797 10192 56831
rect 10140 56788 10192 56797
rect 1492 56695 1544 56704
rect 1492 56661 1501 56695
rect 1501 56661 1535 56695
rect 1535 56661 1544 56695
rect 1492 56652 1544 56661
rect 2228 56695 2280 56704
rect 2228 56661 2237 56695
rect 2237 56661 2271 56695
rect 2271 56661 2280 56695
rect 2228 56652 2280 56661
rect 4213 56550 4265 56602
rect 4277 56550 4329 56602
rect 4341 56550 4393 56602
rect 4405 56550 4457 56602
rect 4469 56550 4521 56602
rect 7477 56550 7529 56602
rect 7541 56550 7593 56602
rect 7605 56550 7657 56602
rect 7669 56550 7721 56602
rect 7733 56550 7785 56602
rect 1400 56448 1452 56500
rect 1676 56448 1728 56500
rect 2596 56423 2648 56432
rect 2596 56389 2605 56423
rect 2605 56389 2639 56423
rect 2639 56389 2648 56423
rect 2596 56380 2648 56389
rect 8852 56448 8904 56500
rect 2964 56380 3016 56432
rect 3608 56380 3660 56432
rect 3240 56312 3292 56364
rect 3516 56355 3568 56364
rect 1400 56244 1452 56296
rect 1952 56244 2004 56296
rect 3516 56321 3525 56355
rect 3525 56321 3559 56355
rect 3559 56321 3568 56355
rect 3516 56312 3568 56321
rect 5264 56244 5316 56296
rect 3240 56176 3292 56228
rect 3884 56176 3936 56228
rect 1400 56108 1452 56160
rect 1952 56108 2004 56160
rect 2136 56108 2188 56160
rect 9864 56108 9916 56160
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5845 56006 5897 56058
rect 5909 56006 5961 56058
rect 5973 56006 6025 56058
rect 6037 56006 6089 56058
rect 6101 56006 6153 56058
rect 9109 56006 9161 56058
rect 9173 56006 9225 56058
rect 9237 56006 9289 56058
rect 9301 56006 9353 56058
rect 9365 56006 9417 56058
rect 2964 55947 3016 55956
rect 2964 55913 2973 55947
rect 2973 55913 3007 55947
rect 3007 55913 3016 55947
rect 2964 55904 3016 55913
rect 4804 55836 4856 55888
rect 8760 55768 8812 55820
rect 3056 55743 3108 55752
rect 3056 55709 3065 55743
rect 3065 55709 3099 55743
rect 3099 55709 3108 55743
rect 3056 55700 3108 55709
rect 10140 55743 10192 55752
rect 10140 55709 10149 55743
rect 10149 55709 10183 55743
rect 10183 55709 10192 55743
rect 10140 55700 10192 55709
rect 1492 55607 1544 55616
rect 1492 55573 1501 55607
rect 1501 55573 1535 55607
rect 1535 55573 1544 55607
rect 1492 55564 1544 55573
rect 2320 55607 2372 55616
rect 2320 55573 2329 55607
rect 2329 55573 2363 55607
rect 2363 55573 2372 55607
rect 2320 55564 2372 55573
rect 4213 55462 4265 55514
rect 4277 55462 4329 55514
rect 4341 55462 4393 55514
rect 4405 55462 4457 55514
rect 4469 55462 4521 55514
rect 7477 55462 7529 55514
rect 7541 55462 7593 55514
rect 7605 55462 7657 55514
rect 7669 55462 7721 55514
rect 7733 55462 7785 55514
rect 1216 55360 1268 55412
rect 1584 55335 1636 55344
rect 1584 55301 1593 55335
rect 1593 55301 1627 55335
rect 1627 55301 1636 55335
rect 1584 55292 1636 55301
rect 3332 55335 3384 55344
rect 3332 55301 3341 55335
rect 3341 55301 3375 55335
rect 3375 55301 3384 55335
rect 3332 55292 3384 55301
rect 2320 55224 2372 55276
rect 3056 55224 3108 55276
rect 1584 55156 1636 55208
rect 10232 55156 10284 55208
rect 2044 55020 2096 55072
rect 9956 55063 10008 55072
rect 9956 55029 9965 55063
rect 9965 55029 9999 55063
rect 9999 55029 10008 55063
rect 9956 55020 10008 55029
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5845 54918 5897 54970
rect 5909 54918 5961 54970
rect 5973 54918 6025 54970
rect 6037 54918 6089 54970
rect 6101 54918 6153 54970
rect 9109 54918 9161 54970
rect 9173 54918 9225 54970
rect 9237 54918 9289 54970
rect 9301 54918 9353 54970
rect 9365 54918 9417 54970
rect 1216 54816 1268 54868
rect 2320 54816 2372 54868
rect 480 54748 532 54800
rect 3608 54748 3660 54800
rect 4712 54612 4764 54664
rect 5448 54544 5500 54596
rect 1400 54476 1452 54528
rect 2780 54476 2832 54528
rect 4213 54374 4265 54426
rect 4277 54374 4329 54426
rect 4341 54374 4393 54426
rect 4405 54374 4457 54426
rect 4469 54374 4521 54426
rect 7477 54374 7529 54426
rect 7541 54374 7593 54426
rect 7605 54374 7657 54426
rect 7669 54374 7721 54426
rect 7733 54374 7785 54426
rect 2872 54136 2924 54188
rect 3516 54136 3568 54188
rect 9864 54179 9916 54188
rect 9864 54145 9873 54179
rect 9873 54145 9907 54179
rect 9907 54145 9916 54179
rect 9864 54136 9916 54145
rect 7104 54068 7156 54120
rect 10048 54043 10100 54052
rect 10048 54009 10057 54043
rect 10057 54009 10091 54043
rect 10091 54009 10100 54043
rect 10048 54000 10100 54009
rect 1492 53975 1544 53984
rect 1492 53941 1501 53975
rect 1501 53941 1535 53975
rect 1535 53941 1544 53975
rect 1492 53932 1544 53941
rect 9864 53932 9916 53984
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5845 53830 5897 53882
rect 5909 53830 5961 53882
rect 5973 53830 6025 53882
rect 6037 53830 6089 53882
rect 6101 53830 6153 53882
rect 9109 53830 9161 53882
rect 9173 53830 9225 53882
rect 9237 53830 9289 53882
rect 9301 53830 9353 53882
rect 9365 53830 9417 53882
rect 1584 53728 1636 53780
rect 1768 53660 1820 53712
rect 1308 53524 1360 53576
rect 1952 53728 2004 53780
rect 8668 53660 8720 53712
rect 3332 53524 3384 53576
rect 1860 53388 1912 53440
rect 2596 53456 2648 53508
rect 2964 53456 3016 53508
rect 9956 53456 10008 53508
rect 10048 53431 10100 53440
rect 10048 53397 10057 53431
rect 10057 53397 10091 53431
rect 10091 53397 10100 53431
rect 10048 53388 10100 53397
rect 4213 53286 4265 53338
rect 4277 53286 4329 53338
rect 4341 53286 4393 53338
rect 4405 53286 4457 53338
rect 4469 53286 4521 53338
rect 7477 53286 7529 53338
rect 7541 53286 7593 53338
rect 7605 53286 7657 53338
rect 7669 53286 7721 53338
rect 7733 53286 7785 53338
rect 7288 53116 7340 53168
rect 1952 53048 2004 53100
rect 7380 53048 7432 53100
rect 9864 53091 9916 53100
rect 9864 53057 9873 53091
rect 9873 53057 9907 53091
rect 9907 53057 9916 53091
rect 9864 53048 9916 53057
rect 296 52912 348 52964
rect 2596 52912 2648 52964
rect 3056 52955 3108 52964
rect 3056 52921 3065 52955
rect 3065 52921 3099 52955
rect 3099 52921 3108 52955
rect 3056 52912 3108 52921
rect 1400 52844 1452 52896
rect 2320 52887 2372 52896
rect 2320 52853 2329 52887
rect 2329 52853 2363 52887
rect 2363 52853 2372 52887
rect 2320 52844 2372 52853
rect 10048 52887 10100 52896
rect 10048 52853 10057 52887
rect 10057 52853 10091 52887
rect 10091 52853 10100 52887
rect 10048 52844 10100 52853
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5845 52742 5897 52794
rect 5909 52742 5961 52794
rect 5973 52742 6025 52794
rect 6037 52742 6089 52794
rect 6101 52742 6153 52794
rect 9109 52742 9161 52794
rect 9173 52742 9225 52794
rect 9237 52742 9289 52794
rect 9301 52742 9353 52794
rect 9365 52742 9417 52794
rect 1952 52640 2004 52692
rect 2228 52683 2280 52692
rect 2228 52649 2237 52683
rect 2237 52649 2271 52683
rect 2271 52649 2280 52683
rect 2228 52640 2280 52649
rect 6276 52572 6328 52624
rect 1860 52436 1912 52488
rect 2596 52504 2648 52556
rect 3332 52504 3384 52556
rect 2320 52436 2372 52488
rect 1492 52343 1544 52352
rect 1492 52309 1501 52343
rect 1501 52309 1535 52343
rect 1535 52309 1544 52343
rect 1492 52300 1544 52309
rect 4213 52198 4265 52250
rect 4277 52198 4329 52250
rect 4341 52198 4393 52250
rect 4405 52198 4457 52250
rect 4469 52198 4521 52250
rect 7477 52198 7529 52250
rect 7541 52198 7593 52250
rect 7605 52198 7657 52250
rect 7669 52198 7721 52250
rect 7733 52198 7785 52250
rect 1768 52096 1820 52148
rect 1952 52096 2004 52148
rect 1308 51960 1360 52012
rect 2596 52003 2648 52012
rect 1584 51824 1636 51876
rect 2596 51969 2605 52003
rect 2605 51969 2639 52003
rect 2639 51969 2648 52003
rect 2596 51960 2648 51969
rect 2964 51960 3016 52012
rect 3516 51960 3568 52012
rect 480 51756 532 51808
rect 3332 51824 3384 51876
rect 10048 51799 10100 51808
rect 10048 51765 10057 51799
rect 10057 51765 10091 51799
rect 10091 51765 10100 51799
rect 10048 51756 10100 51765
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5845 51654 5897 51706
rect 5909 51654 5961 51706
rect 5973 51654 6025 51706
rect 6037 51654 6089 51706
rect 6101 51654 6153 51706
rect 9109 51654 9161 51706
rect 9173 51654 9225 51706
rect 9237 51654 9289 51706
rect 9301 51654 9353 51706
rect 9365 51654 9417 51706
rect 7932 51416 7984 51468
rect 2780 51348 2832 51400
rect 9864 51391 9916 51400
rect 9864 51357 9873 51391
rect 9873 51357 9907 51391
rect 9907 51357 9916 51391
rect 9864 51348 9916 51357
rect 7840 51280 7892 51332
rect 1400 51212 1452 51264
rect 2228 51255 2280 51264
rect 2228 51221 2237 51255
rect 2237 51221 2271 51255
rect 2271 51221 2280 51255
rect 2228 51212 2280 51221
rect 3056 51255 3108 51264
rect 3056 51221 3065 51255
rect 3065 51221 3099 51255
rect 3099 51221 3108 51255
rect 3056 51212 3108 51221
rect 10048 51255 10100 51264
rect 10048 51221 10057 51255
rect 10057 51221 10091 51255
rect 10091 51221 10100 51255
rect 10048 51212 10100 51221
rect 4213 51110 4265 51162
rect 4277 51110 4329 51162
rect 4341 51110 4393 51162
rect 4405 51110 4457 51162
rect 4469 51110 4521 51162
rect 7477 51110 7529 51162
rect 7541 51110 7593 51162
rect 7605 51110 7657 51162
rect 7669 51110 7721 51162
rect 7733 51110 7785 51162
rect 9864 51008 9916 51060
rect 3516 50940 3568 50992
rect 4160 50872 4212 50924
rect 7196 50804 7248 50856
rect 2780 50736 2832 50788
rect 3792 50736 3844 50788
rect 1492 50711 1544 50720
rect 1492 50677 1501 50711
rect 1501 50677 1535 50711
rect 1535 50677 1544 50711
rect 1492 50668 1544 50677
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5845 50566 5897 50618
rect 5909 50566 5961 50618
rect 5973 50566 6025 50618
rect 6037 50566 6089 50618
rect 6101 50566 6153 50618
rect 9109 50566 9161 50618
rect 9173 50566 9225 50618
rect 9237 50566 9289 50618
rect 9301 50566 9353 50618
rect 9365 50566 9417 50618
rect 1308 50464 1360 50516
rect 1952 50464 2004 50516
rect 2504 50464 2556 50516
rect 3700 50464 3752 50516
rect 1676 50396 1728 50448
rect 2412 50396 2464 50448
rect 3516 50396 3568 50448
rect 1308 50328 1360 50380
rect 1584 50303 1636 50312
rect 1584 50269 1593 50303
rect 1593 50269 1627 50303
rect 1627 50269 1636 50303
rect 1584 50260 1636 50269
rect 1032 50192 1084 50244
rect 1952 50303 2004 50312
rect 1952 50269 1961 50303
rect 1961 50269 1995 50303
rect 1995 50269 2004 50303
rect 1952 50260 2004 50269
rect 2964 50260 3016 50312
rect 1676 50124 1728 50176
rect 4160 50192 4212 50244
rect 4620 50192 4672 50244
rect 10048 50167 10100 50176
rect 10048 50133 10057 50167
rect 10057 50133 10091 50167
rect 10091 50133 10100 50167
rect 10048 50124 10100 50133
rect 4213 50022 4265 50074
rect 4277 50022 4329 50074
rect 4341 50022 4393 50074
rect 4405 50022 4457 50074
rect 4469 50022 4521 50074
rect 7477 50022 7529 50074
rect 7541 50022 7593 50074
rect 7605 50022 7657 50074
rect 7669 50022 7721 50074
rect 7733 50022 7785 50074
rect 1584 49827 1636 49836
rect 1584 49793 1593 49827
rect 1593 49793 1627 49827
rect 1627 49793 1636 49827
rect 1584 49784 1636 49793
rect 1952 49827 2004 49836
rect 1124 49716 1176 49768
rect 1952 49793 1961 49827
rect 1961 49793 1995 49827
rect 1995 49793 2004 49827
rect 1952 49784 2004 49793
rect 6184 49784 6236 49836
rect 9864 49827 9916 49836
rect 9864 49793 9873 49827
rect 9873 49793 9907 49827
rect 9907 49793 9916 49827
rect 9864 49784 9916 49793
rect 1492 49648 1544 49700
rect 3976 49716 4028 49768
rect 5172 49716 5224 49768
rect 1400 49623 1452 49632
rect 1400 49589 1409 49623
rect 1409 49589 1443 49623
rect 1443 49589 1452 49623
rect 1400 49580 1452 49589
rect 1952 49580 2004 49632
rect 2320 49580 2372 49632
rect 2412 49580 2464 49632
rect 4620 49580 4672 49632
rect 5172 49580 5224 49632
rect 10048 49623 10100 49632
rect 10048 49589 10057 49623
rect 10057 49589 10091 49623
rect 10091 49589 10100 49623
rect 10048 49580 10100 49589
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5845 49478 5897 49530
rect 5909 49478 5961 49530
rect 5973 49478 6025 49530
rect 6037 49478 6089 49530
rect 6101 49478 6153 49530
rect 9109 49478 9161 49530
rect 9173 49478 9225 49530
rect 9237 49478 9289 49530
rect 9301 49478 9353 49530
rect 9365 49478 9417 49530
rect 1492 49172 1544 49224
rect 6736 49240 6788 49292
rect 388 49104 440 49156
rect 3516 49172 3568 49224
rect 4620 49172 4672 49224
rect 9772 49172 9824 49224
rect 1492 49036 1544 49088
rect 2320 49036 2372 49088
rect 2780 49036 2832 49088
rect 3516 49036 3568 49088
rect 10048 49079 10100 49088
rect 10048 49045 10057 49079
rect 10057 49045 10091 49079
rect 10091 49045 10100 49079
rect 10048 49036 10100 49045
rect 4213 48934 4265 48986
rect 4277 48934 4329 48986
rect 4341 48934 4393 48986
rect 4405 48934 4457 48986
rect 4469 48934 4521 48986
rect 7477 48934 7529 48986
rect 7541 48934 7593 48986
rect 7605 48934 7657 48986
rect 7669 48934 7721 48986
rect 7733 48934 7785 48986
rect 388 48832 440 48884
rect 1308 48832 1360 48884
rect 2228 48875 2280 48884
rect 2228 48841 2237 48875
rect 2237 48841 2271 48875
rect 2271 48841 2280 48875
rect 2228 48832 2280 48841
rect 6552 48696 6604 48748
rect 6460 48628 6512 48680
rect 2228 48560 2280 48612
rect 2412 48560 2464 48612
rect 1492 48535 1544 48544
rect 1492 48501 1501 48535
rect 1501 48501 1535 48535
rect 1535 48501 1544 48535
rect 1492 48492 1544 48501
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5845 48390 5897 48442
rect 5909 48390 5961 48442
rect 5973 48390 6025 48442
rect 6037 48390 6089 48442
rect 6101 48390 6153 48442
rect 9109 48390 9161 48442
rect 9173 48390 9225 48442
rect 9237 48390 9289 48442
rect 9301 48390 9353 48442
rect 9365 48390 9417 48442
rect 20 48288 72 48340
rect 1584 48288 1636 48340
rect 2412 48288 2464 48340
rect 5540 48288 5592 48340
rect 2872 48220 2924 48272
rect 3056 48220 3108 48272
rect 4528 48152 4580 48204
rect 1952 48084 2004 48136
rect 2780 48127 2832 48136
rect 2780 48093 2789 48127
rect 2789 48093 2823 48127
rect 2823 48093 2832 48127
rect 2780 48084 2832 48093
rect 3056 48084 3108 48136
rect 6184 48016 6236 48068
rect 1492 47991 1544 48000
rect 1492 47957 1501 47991
rect 1501 47957 1535 47991
rect 1535 47957 1544 47991
rect 1492 47948 1544 47957
rect 9864 47948 9916 48000
rect 10048 47991 10100 48000
rect 10048 47957 10057 47991
rect 10057 47957 10091 47991
rect 10091 47957 10100 47991
rect 10048 47948 10100 47957
rect 4213 47846 4265 47898
rect 4277 47846 4329 47898
rect 4341 47846 4393 47898
rect 4405 47846 4457 47898
rect 4469 47846 4521 47898
rect 7477 47846 7529 47898
rect 7541 47846 7593 47898
rect 7605 47846 7657 47898
rect 7669 47846 7721 47898
rect 7733 47846 7785 47898
rect 2964 47787 3016 47796
rect 2964 47753 2973 47787
rect 2973 47753 3007 47787
rect 3007 47753 3016 47787
rect 2964 47744 3016 47753
rect 3516 47744 3568 47796
rect 2504 47676 2556 47728
rect 1308 47608 1360 47660
rect 2688 47608 2740 47660
rect 2872 47651 2924 47660
rect 2872 47617 2881 47651
rect 2881 47617 2915 47651
rect 2915 47617 2924 47651
rect 2872 47608 2924 47617
rect 2964 47608 3016 47660
rect 3516 47651 3568 47660
rect 3516 47617 3525 47651
rect 3525 47617 3559 47651
rect 3559 47617 3568 47651
rect 3516 47608 3568 47617
rect 1492 47540 1544 47592
rect 2136 47472 2188 47524
rect 2504 47540 2556 47592
rect 1492 47447 1544 47456
rect 1492 47413 1501 47447
rect 1501 47413 1535 47447
rect 1535 47413 1544 47447
rect 1492 47404 1544 47413
rect 10048 47447 10100 47456
rect 10048 47413 10057 47447
rect 10057 47413 10091 47447
rect 10091 47413 10100 47447
rect 10048 47404 10100 47413
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5845 47302 5897 47354
rect 5909 47302 5961 47354
rect 5973 47302 6025 47354
rect 6037 47302 6089 47354
rect 6101 47302 6153 47354
rect 9109 47302 9161 47354
rect 9173 47302 9225 47354
rect 9237 47302 9289 47354
rect 9301 47302 9353 47354
rect 9365 47302 9417 47354
rect 3056 47243 3108 47252
rect 3056 47209 3065 47243
rect 3065 47209 3099 47243
rect 3099 47209 3108 47243
rect 3056 47200 3108 47209
rect 1952 47132 2004 47184
rect 2228 47132 2280 47184
rect 1032 47064 1084 47116
rect 3516 47132 3568 47184
rect 1492 46903 1544 46912
rect 1492 46869 1501 46903
rect 1501 46869 1535 46903
rect 1535 46869 1544 46903
rect 1492 46860 1544 46869
rect 2504 46996 2556 47048
rect 2872 47039 2924 47048
rect 2872 47005 2881 47039
rect 2881 47005 2915 47039
rect 2915 47005 2924 47039
rect 2872 46996 2924 47005
rect 2596 46860 2648 46912
rect 2780 46860 2832 46912
rect 4213 46758 4265 46810
rect 4277 46758 4329 46810
rect 4341 46758 4393 46810
rect 4405 46758 4457 46810
rect 4469 46758 4521 46810
rect 7477 46758 7529 46810
rect 7541 46758 7593 46810
rect 7605 46758 7657 46810
rect 7669 46758 7721 46810
rect 7733 46758 7785 46810
rect 1124 46656 1176 46708
rect 2872 46656 2924 46708
rect 2596 46588 2648 46640
rect 8944 46588 8996 46640
rect 1952 46520 2004 46572
rect 2780 46520 2832 46572
rect 3516 46520 3568 46572
rect 3792 46520 3844 46572
rect 9036 46452 9088 46504
rect 9772 46384 9824 46436
rect 10048 46427 10100 46436
rect 10048 46393 10057 46427
rect 10057 46393 10091 46427
rect 10091 46393 10100 46427
rect 10048 46384 10100 46393
rect 1492 46359 1544 46368
rect 1492 46325 1501 46359
rect 1501 46325 1535 46359
rect 1535 46325 1544 46359
rect 1492 46316 1544 46325
rect 4620 46316 4672 46368
rect 5356 46316 5408 46368
rect 388 46248 440 46300
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5845 46214 5897 46266
rect 5909 46214 5961 46266
rect 5973 46214 6025 46266
rect 6037 46214 6089 46266
rect 6101 46214 6153 46266
rect 9109 46214 9161 46266
rect 9173 46214 9225 46266
rect 9237 46214 9289 46266
rect 9301 46214 9353 46266
rect 9365 46214 9417 46266
rect 4804 46112 4856 46164
rect 4988 46112 5040 46164
rect 112 46044 164 46096
rect 480 46044 532 46096
rect 1216 46044 1268 46096
rect 3608 46044 3660 46096
rect 4068 46044 4120 46096
rect 4528 46044 4580 46096
rect 5356 46044 5408 46096
rect 4712 45976 4764 46028
rect 4988 45976 5040 46028
rect 8024 45908 8076 45960
rect 9864 45951 9916 45960
rect 9864 45917 9873 45951
rect 9873 45917 9907 45951
rect 9907 45917 9916 45951
rect 9864 45908 9916 45917
rect 4712 45840 4764 45892
rect 5448 45840 5500 45892
rect 1492 45815 1544 45824
rect 1492 45781 1501 45815
rect 1501 45781 1535 45815
rect 1535 45781 1544 45815
rect 1492 45772 1544 45781
rect 10048 45815 10100 45824
rect 10048 45781 10057 45815
rect 10057 45781 10091 45815
rect 10091 45781 10100 45815
rect 10048 45772 10100 45781
rect 4213 45670 4265 45722
rect 4277 45670 4329 45722
rect 4341 45670 4393 45722
rect 4405 45670 4457 45722
rect 4469 45670 4521 45722
rect 7477 45670 7529 45722
rect 7541 45670 7593 45722
rect 7605 45670 7657 45722
rect 7669 45670 7721 45722
rect 7733 45670 7785 45722
rect 1676 45568 1728 45620
rect 1952 45568 2004 45620
rect 5172 45568 5224 45620
rect 5356 45568 5408 45620
rect 3424 45500 3476 45552
rect 1952 45432 2004 45484
rect 1492 45271 1544 45280
rect 1492 45237 1501 45271
rect 1501 45237 1535 45271
rect 1535 45237 1544 45271
rect 1492 45228 1544 45237
rect 1860 45228 1912 45280
rect 5632 45228 5684 45280
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5845 45126 5897 45178
rect 5909 45126 5961 45178
rect 5973 45126 6025 45178
rect 6037 45126 6089 45178
rect 6101 45126 6153 45178
rect 9109 45126 9161 45178
rect 9173 45126 9225 45178
rect 9237 45126 9289 45178
rect 9301 45126 9353 45178
rect 9365 45126 9417 45178
rect 1492 45024 1544 45076
rect 4068 45024 4120 45076
rect 5080 45024 5132 45076
rect 1768 44956 1820 45008
rect 2504 44956 2556 45008
rect 2780 44956 2832 45008
rect 2228 44888 2280 44940
rect 6828 44820 6880 44872
rect 9680 44820 9732 44872
rect 2780 44684 2832 44736
rect 10048 44727 10100 44736
rect 10048 44693 10057 44727
rect 10057 44693 10091 44727
rect 10091 44693 10100 44727
rect 10048 44684 10100 44693
rect 4213 44582 4265 44634
rect 4277 44582 4329 44634
rect 4341 44582 4393 44634
rect 4405 44582 4457 44634
rect 4469 44582 4521 44634
rect 7477 44582 7529 44634
rect 7541 44582 7593 44634
rect 7605 44582 7657 44634
rect 7669 44582 7721 44634
rect 7733 44582 7785 44634
rect 1492 44523 1544 44532
rect 1492 44489 1501 44523
rect 1501 44489 1535 44523
rect 1535 44489 1544 44523
rect 1492 44480 1544 44489
rect 1768 44344 1820 44396
rect 2412 44344 2464 44396
rect 3148 44387 3200 44396
rect 3148 44353 3157 44387
rect 3157 44353 3191 44387
rect 3191 44353 3200 44387
rect 3148 44344 3200 44353
rect 4160 44344 4212 44396
rect 9772 44344 9824 44396
rect 9680 44276 9732 44328
rect 2136 44208 2188 44260
rect 2412 44208 2464 44260
rect 5540 44208 5592 44260
rect 2320 44183 2372 44192
rect 2320 44149 2329 44183
rect 2329 44149 2363 44183
rect 2363 44149 2372 44183
rect 2320 44140 2372 44149
rect 2964 44183 3016 44192
rect 2964 44149 2973 44183
rect 2973 44149 3007 44183
rect 3007 44149 3016 44183
rect 2964 44140 3016 44149
rect 3240 44140 3292 44192
rect 3792 44140 3844 44192
rect 10048 44183 10100 44192
rect 10048 44149 10057 44183
rect 10057 44149 10091 44183
rect 10091 44149 10100 44183
rect 10048 44140 10100 44149
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5845 44038 5897 44090
rect 5909 44038 5961 44090
rect 5973 44038 6025 44090
rect 6037 44038 6089 44090
rect 6101 44038 6153 44090
rect 9109 44038 9161 44090
rect 9173 44038 9225 44090
rect 9237 44038 9289 44090
rect 9301 44038 9353 44090
rect 9365 44038 9417 44090
rect 572 43936 624 43988
rect 1216 43936 1268 43988
rect 5540 43936 5592 43988
rect 6184 43936 6236 43988
rect 2136 43800 2188 43852
rect 2504 43800 2556 43852
rect 6184 43800 6236 43852
rect 6736 43800 6788 43852
rect 1676 43732 1728 43784
rect 1860 43732 1912 43784
rect 572 43664 624 43716
rect 3608 43732 3660 43784
rect 4160 43732 4212 43784
rect 9588 43732 9640 43784
rect 2964 43664 3016 43716
rect 8300 43664 8352 43716
rect 2780 43596 2832 43648
rect 9680 43596 9732 43648
rect 10048 43639 10100 43648
rect 10048 43605 10057 43639
rect 10057 43605 10091 43639
rect 10091 43605 10100 43639
rect 10048 43596 10100 43605
rect 4213 43494 4265 43546
rect 4277 43494 4329 43546
rect 4341 43494 4393 43546
rect 4405 43494 4457 43546
rect 4469 43494 4521 43546
rect 7477 43494 7529 43546
rect 7541 43494 7593 43546
rect 7605 43494 7657 43546
rect 7669 43494 7721 43546
rect 7733 43494 7785 43546
rect 3884 43392 3936 43444
rect 9864 43392 9916 43444
rect 940 43324 992 43376
rect 2136 43324 2188 43376
rect 940 43188 992 43240
rect 1124 43188 1176 43240
rect 2964 43324 3016 43376
rect 3056 43324 3108 43376
rect 9772 43324 9824 43376
rect 572 43120 624 43172
rect 3608 43256 3660 43308
rect 3884 43299 3936 43308
rect 3884 43265 3893 43299
rect 3893 43265 3927 43299
rect 3927 43265 3936 43299
rect 3884 43256 3936 43265
rect 4160 43256 4212 43308
rect 3608 43120 3660 43172
rect 2964 43052 3016 43104
rect 4160 43052 4212 43104
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5845 42950 5897 43002
rect 5909 42950 5961 43002
rect 5973 42950 6025 43002
rect 6037 42950 6089 43002
rect 6101 42950 6153 43002
rect 9109 42950 9161 43002
rect 9173 42950 9225 43002
rect 9237 42950 9289 43002
rect 9301 42950 9353 43002
rect 9365 42950 9417 43002
rect 2872 42780 2924 42832
rect 2136 42687 2188 42696
rect 2136 42653 2145 42687
rect 2145 42653 2179 42687
rect 2179 42653 2188 42687
rect 2136 42644 2188 42653
rect 1676 42576 1728 42628
rect 3700 42644 3752 42696
rect 4160 42848 4212 42900
rect 9680 42780 9732 42832
rect 2504 42576 2556 42628
rect 848 42508 900 42560
rect 3056 42551 3108 42560
rect 3056 42517 3065 42551
rect 3065 42517 3099 42551
rect 3099 42517 3108 42551
rect 3056 42508 3108 42517
rect 10048 42551 10100 42560
rect 10048 42517 10057 42551
rect 10057 42517 10091 42551
rect 10091 42517 10100 42551
rect 10048 42508 10100 42517
rect 4213 42406 4265 42458
rect 4277 42406 4329 42458
rect 4341 42406 4393 42458
rect 4405 42406 4457 42458
rect 4469 42406 4521 42458
rect 7477 42406 7529 42458
rect 7541 42406 7593 42458
rect 7605 42406 7657 42458
rect 7669 42406 7721 42458
rect 7733 42406 7785 42458
rect 9588 42304 9640 42356
rect 2412 42211 2464 42220
rect 2412 42177 2421 42211
rect 2421 42177 2455 42211
rect 2455 42177 2464 42211
rect 2412 42168 2464 42177
rect 2964 42236 3016 42288
rect 9864 42211 9916 42220
rect 9864 42177 9873 42211
rect 9873 42177 9907 42211
rect 9907 42177 9916 42211
rect 9864 42168 9916 42177
rect 1676 42032 1728 42084
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 2228 42007 2280 42016
rect 2228 41973 2237 42007
rect 2237 41973 2271 42007
rect 2271 41973 2280 42007
rect 2228 41964 2280 41973
rect 10048 42007 10100 42016
rect 10048 41973 10057 42007
rect 10057 41973 10091 42007
rect 10091 41973 10100 42007
rect 10048 41964 10100 41973
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5845 41862 5897 41914
rect 5909 41862 5961 41914
rect 5973 41862 6025 41914
rect 6037 41862 6089 41914
rect 6101 41862 6153 41914
rect 9109 41862 9161 41914
rect 9173 41862 9225 41914
rect 9237 41862 9289 41914
rect 9301 41862 9353 41914
rect 9365 41862 9417 41914
rect 9864 41760 9916 41812
rect 1860 41692 1912 41744
rect 3792 41692 3844 41744
rect 204 41624 256 41676
rect 2228 41624 2280 41676
rect 1768 41556 1820 41608
rect 1860 41556 1912 41608
rect 2136 41599 2188 41608
rect 204 41531 256 41540
rect 204 41497 213 41531
rect 213 41497 247 41531
rect 247 41497 256 41531
rect 204 41488 256 41497
rect 2136 41565 2145 41599
rect 2145 41565 2179 41599
rect 2179 41565 2188 41599
rect 2136 41556 2188 41565
rect 2688 41624 2740 41676
rect 7012 41624 7064 41676
rect 2964 41599 3016 41608
rect 2964 41565 2973 41599
rect 2973 41565 3007 41599
rect 3007 41565 3016 41599
rect 2964 41556 3016 41565
rect 1216 41420 1268 41472
rect 1768 41420 1820 41472
rect 3608 41488 3660 41540
rect 2412 41420 2464 41472
rect 3424 41420 3476 41472
rect 5724 41420 5776 41472
rect 4213 41318 4265 41370
rect 4277 41318 4329 41370
rect 4341 41318 4393 41370
rect 4405 41318 4457 41370
rect 4469 41318 4521 41370
rect 7477 41318 7529 41370
rect 7541 41318 7593 41370
rect 7605 41318 7657 41370
rect 7669 41318 7721 41370
rect 7733 41318 7785 41370
rect 3332 41216 3384 41268
rect 3976 41216 4028 41268
rect 8392 41148 8444 41200
rect 2688 41080 2740 41132
rect 4068 41080 4120 41132
rect 9680 41080 9732 41132
rect 2044 41012 2096 41064
rect 2228 41012 2280 41064
rect 3056 40987 3108 40996
rect 3056 40953 3065 40987
rect 3065 40953 3099 40987
rect 3099 40953 3108 40987
rect 3056 40944 3108 40953
rect 10048 40987 10100 40996
rect 10048 40953 10057 40987
rect 10057 40953 10091 40987
rect 10091 40953 10100 40987
rect 10048 40944 10100 40953
rect 1216 40876 1268 40928
rect 2228 40919 2280 40928
rect 2228 40885 2237 40919
rect 2237 40885 2271 40919
rect 2271 40885 2280 40919
rect 2228 40876 2280 40885
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5845 40774 5897 40826
rect 5909 40774 5961 40826
rect 5973 40774 6025 40826
rect 6037 40774 6089 40826
rect 6101 40774 6153 40826
rect 9109 40774 9161 40826
rect 9173 40774 9225 40826
rect 9237 40774 9289 40826
rect 9301 40774 9353 40826
rect 9365 40774 9417 40826
rect 664 40672 716 40724
rect 1768 40468 1820 40520
rect 2872 40468 2924 40520
rect 9864 40511 9916 40520
rect 9864 40477 9873 40511
rect 9873 40477 9907 40511
rect 9907 40477 9916 40511
rect 9864 40468 9916 40477
rect 2596 40400 2648 40452
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 10048 40375 10100 40384
rect 10048 40341 10057 40375
rect 10057 40341 10091 40375
rect 10091 40341 10100 40375
rect 10048 40332 10100 40341
rect 4213 40230 4265 40282
rect 4277 40230 4329 40282
rect 4341 40230 4393 40282
rect 4405 40230 4457 40282
rect 4469 40230 4521 40282
rect 7477 40230 7529 40282
rect 7541 40230 7593 40282
rect 7605 40230 7657 40282
rect 7669 40230 7721 40282
rect 7733 40230 7785 40282
rect 1860 40128 1912 40180
rect 2596 40128 2648 40180
rect 4804 40060 4856 40112
rect 1860 39992 1912 40044
rect 2320 40035 2372 40044
rect 2320 40001 2329 40035
rect 2329 40001 2363 40035
rect 2363 40001 2372 40035
rect 2872 40035 2924 40044
rect 2320 39992 2372 40001
rect 2872 40001 2881 40035
rect 2881 40001 2915 40035
rect 2915 40001 2924 40035
rect 2872 39992 2924 40001
rect 3056 40035 3108 40044
rect 3056 40001 3065 40035
rect 3065 40001 3099 40035
rect 3099 40001 3108 40035
rect 3056 39992 3108 40001
rect 9772 39992 9824 40044
rect 1216 39788 1268 39840
rect 9680 39856 9732 39908
rect 2228 39788 2280 39840
rect 10048 39831 10100 39840
rect 10048 39797 10057 39831
rect 10057 39797 10091 39831
rect 10091 39797 10100 39831
rect 10048 39788 10100 39797
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5845 39686 5897 39738
rect 5909 39686 5961 39738
rect 5973 39686 6025 39738
rect 6037 39686 6089 39738
rect 6101 39686 6153 39738
rect 9109 39686 9161 39738
rect 9173 39686 9225 39738
rect 9237 39686 9289 39738
rect 9301 39686 9353 39738
rect 9365 39686 9417 39738
rect 20 39448 72 39500
rect 1492 39380 1544 39432
rect 1860 39380 1912 39432
rect 3424 39380 3476 39432
rect 2872 39312 2924 39364
rect 2780 39244 2832 39296
rect 4213 39142 4265 39194
rect 4277 39142 4329 39194
rect 4341 39142 4393 39194
rect 4405 39142 4457 39194
rect 4469 39142 4521 39194
rect 7477 39142 7529 39194
rect 7541 39142 7593 39194
rect 7605 39142 7657 39194
rect 7669 39142 7721 39194
rect 7733 39142 7785 39194
rect 3516 39040 3568 39092
rect 9864 39040 9916 39092
rect 1860 38947 1912 38956
rect 1860 38913 1869 38947
rect 1869 38913 1903 38947
rect 1903 38913 1912 38947
rect 1860 38904 1912 38913
rect 3608 38972 3660 39024
rect 3240 38947 3292 38956
rect 3240 38913 3249 38947
rect 3249 38913 3283 38947
rect 3283 38913 3292 38947
rect 3240 38904 3292 38913
rect 2964 38836 3016 38888
rect 3516 38836 3568 38888
rect 2872 38768 2924 38820
rect 3240 38768 3292 38820
rect 4068 38904 4120 38956
rect 9864 38947 9916 38956
rect 9864 38913 9873 38947
rect 9873 38913 9907 38947
rect 9907 38913 9916 38947
rect 9864 38904 9916 38913
rect 2964 38700 3016 38752
rect 3424 38743 3476 38752
rect 3424 38709 3433 38743
rect 3433 38709 3467 38743
rect 3467 38709 3476 38743
rect 3424 38700 3476 38709
rect 3700 38700 3752 38752
rect 6368 38700 6420 38752
rect 10048 38743 10100 38752
rect 10048 38709 10057 38743
rect 10057 38709 10091 38743
rect 10091 38709 10100 38743
rect 10048 38700 10100 38709
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5845 38598 5897 38650
rect 5909 38598 5961 38650
rect 5973 38598 6025 38650
rect 6037 38598 6089 38650
rect 6101 38598 6153 38650
rect 9109 38598 9161 38650
rect 9173 38598 9225 38650
rect 9237 38598 9289 38650
rect 9301 38598 9353 38650
rect 9365 38598 9417 38650
rect 1124 38496 1176 38548
rect 1492 38360 1544 38412
rect 2136 38403 2188 38412
rect 1492 38199 1544 38208
rect 1492 38165 1501 38199
rect 1501 38165 1535 38199
rect 1535 38165 1544 38199
rect 1492 38156 1544 38165
rect 2136 38369 2145 38403
rect 2145 38369 2179 38403
rect 2179 38369 2188 38403
rect 2136 38360 2188 38369
rect 9772 38496 9824 38548
rect 2136 38224 2188 38276
rect 3056 38292 3108 38344
rect 3608 38292 3660 38344
rect 4068 38292 4120 38344
rect 3424 38156 3476 38208
rect 10048 38199 10100 38208
rect 10048 38165 10057 38199
rect 10057 38165 10091 38199
rect 10091 38165 10100 38199
rect 10048 38156 10100 38165
rect 4213 38054 4265 38106
rect 4277 38054 4329 38106
rect 4341 38054 4393 38106
rect 4405 38054 4457 38106
rect 4469 38054 4521 38106
rect 7477 38054 7529 38106
rect 7541 38054 7593 38106
rect 7605 38054 7657 38106
rect 7669 38054 7721 38106
rect 7733 38054 7785 38106
rect 756 37952 808 38004
rect 4896 37952 4948 38004
rect 2136 37816 2188 37868
rect 2964 37816 3016 37868
rect 3424 37816 3476 37868
rect 3608 37748 3660 37800
rect 1492 37655 1544 37664
rect 1492 37621 1501 37655
rect 1501 37621 1535 37655
rect 1535 37621 1544 37655
rect 1492 37612 1544 37621
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5845 37510 5897 37562
rect 5909 37510 5961 37562
rect 5973 37510 6025 37562
rect 6037 37510 6089 37562
rect 6101 37510 6153 37562
rect 9109 37510 9161 37562
rect 9173 37510 9225 37562
rect 9237 37510 9289 37562
rect 9301 37510 9353 37562
rect 9365 37510 9417 37562
rect 1032 37204 1084 37256
rect 2136 37340 2188 37392
rect 2964 37340 3016 37392
rect 9864 37340 9916 37392
rect 3056 37204 3108 37256
rect 3240 37204 3292 37256
rect 4620 37136 4672 37188
rect 10048 37111 10100 37120
rect 10048 37077 10057 37111
rect 10057 37077 10091 37111
rect 10091 37077 10100 37111
rect 10048 37068 10100 37077
rect 4213 36966 4265 37018
rect 4277 36966 4329 37018
rect 4341 36966 4393 37018
rect 4405 36966 4457 37018
rect 4469 36966 4521 37018
rect 7477 36966 7529 37018
rect 7541 36966 7593 37018
rect 7605 36966 7657 37018
rect 7669 36966 7721 37018
rect 7733 36966 7785 37018
rect 2320 36796 2372 36848
rect 6920 36796 6972 36848
rect 572 36660 624 36712
rect 1216 36660 1268 36712
rect 9772 36728 9824 36780
rect 8484 36660 8536 36712
rect 3056 36635 3108 36644
rect 3056 36601 3065 36635
rect 3065 36601 3099 36635
rect 3099 36601 3108 36635
rect 3056 36592 3108 36601
rect 204 36524 256 36576
rect 572 36524 624 36576
rect 1492 36567 1544 36576
rect 1492 36533 1501 36567
rect 1501 36533 1535 36567
rect 1535 36533 1544 36567
rect 1492 36524 1544 36533
rect 2320 36567 2372 36576
rect 2320 36533 2329 36567
rect 2329 36533 2363 36567
rect 2363 36533 2372 36567
rect 2320 36524 2372 36533
rect 10048 36567 10100 36576
rect 10048 36533 10057 36567
rect 10057 36533 10091 36567
rect 10091 36533 10100 36567
rect 10048 36524 10100 36533
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5845 36422 5897 36474
rect 5909 36422 5961 36474
rect 5973 36422 6025 36474
rect 6037 36422 6089 36474
rect 6101 36422 6153 36474
rect 9109 36422 9161 36474
rect 9173 36422 9225 36474
rect 9237 36422 9289 36474
rect 9301 36422 9353 36474
rect 9365 36422 9417 36474
rect 3240 36363 3292 36372
rect 3240 36329 3249 36363
rect 3249 36329 3283 36363
rect 3283 36329 3292 36363
rect 3240 36320 3292 36329
rect 4988 36252 5040 36304
rect 756 36184 808 36236
rect 1124 36184 1176 36236
rect 3976 36116 4028 36168
rect 9864 36159 9916 36168
rect 9864 36125 9873 36159
rect 9873 36125 9907 36159
rect 9907 36125 9916 36159
rect 9864 36116 9916 36125
rect 3608 36048 3660 36100
rect 2964 35980 3016 36032
rect 10048 36023 10100 36032
rect 10048 35989 10057 36023
rect 10057 35989 10091 36023
rect 10091 35989 10100 36023
rect 10048 35980 10100 35989
rect 4213 35878 4265 35930
rect 4277 35878 4329 35930
rect 4341 35878 4393 35930
rect 4405 35878 4457 35930
rect 4469 35878 4521 35930
rect 7477 35878 7529 35930
rect 7541 35878 7593 35930
rect 7605 35878 7657 35930
rect 7669 35878 7721 35930
rect 7733 35878 7785 35930
rect 4712 35776 4764 35828
rect 2320 35683 2372 35692
rect 2320 35649 2329 35683
rect 2329 35649 2363 35683
rect 2363 35649 2372 35683
rect 2320 35640 2372 35649
rect 3700 35640 3752 35692
rect 2964 35572 3016 35624
rect 3056 35547 3108 35556
rect 3056 35513 3065 35547
rect 3065 35513 3099 35547
rect 3099 35513 3108 35547
rect 3056 35504 3108 35513
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5845 35334 5897 35386
rect 5909 35334 5961 35386
rect 5973 35334 6025 35386
rect 6037 35334 6089 35386
rect 6101 35334 6153 35386
rect 9109 35334 9161 35386
rect 9173 35334 9225 35386
rect 9237 35334 9289 35386
rect 9301 35334 9353 35386
rect 9365 35334 9417 35386
rect 9864 35232 9916 35284
rect 8852 35164 8904 35216
rect 2136 35071 2188 35080
rect 2136 35037 2145 35071
rect 2145 35037 2179 35071
rect 2179 35037 2188 35071
rect 2136 35028 2188 35037
rect 2964 35028 3016 35080
rect 3608 35028 3660 35080
rect 3976 35071 4028 35080
rect 3976 35037 3985 35071
rect 3985 35037 4019 35071
rect 4019 35037 4028 35071
rect 3976 35028 4028 35037
rect 9864 35071 9916 35080
rect 9864 35037 9873 35071
rect 9873 35037 9907 35071
rect 9907 35037 9916 35071
rect 9864 35028 9916 35037
rect 5448 34960 5500 35012
rect 2964 34892 3016 34944
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 4213 34790 4265 34842
rect 4277 34790 4329 34842
rect 4341 34790 4393 34842
rect 4405 34790 4457 34842
rect 4469 34790 4521 34842
rect 7477 34790 7529 34842
rect 7541 34790 7593 34842
rect 7605 34790 7657 34842
rect 7669 34790 7721 34842
rect 7733 34790 7785 34842
rect 3056 34688 3108 34740
rect 3240 34731 3292 34740
rect 3240 34697 3249 34731
rect 3249 34697 3283 34731
rect 3283 34697 3292 34731
rect 3240 34688 3292 34697
rect 8760 34620 8812 34672
rect 2136 34552 2188 34604
rect 2412 34552 2464 34604
rect 3148 34552 3200 34604
rect 9680 34552 9732 34604
rect 2136 34416 2188 34468
rect 2412 34391 2464 34400
rect 2412 34357 2421 34391
rect 2421 34357 2455 34391
rect 2455 34357 2464 34391
rect 2412 34348 2464 34357
rect 10048 34391 10100 34400
rect 10048 34357 10057 34391
rect 10057 34357 10091 34391
rect 10091 34357 10100 34391
rect 10048 34348 10100 34357
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5845 34246 5897 34298
rect 5909 34246 5961 34298
rect 5973 34246 6025 34298
rect 6037 34246 6089 34298
rect 6101 34246 6153 34298
rect 9109 34246 9161 34298
rect 9173 34246 9225 34298
rect 9237 34246 9289 34298
rect 9301 34246 9353 34298
rect 9365 34246 9417 34298
rect 1492 34187 1544 34196
rect 1492 34153 1501 34187
rect 1501 34153 1535 34187
rect 1535 34153 1544 34187
rect 1492 34144 1544 34153
rect 9772 34144 9824 34196
rect 8576 34076 8628 34128
rect 2136 33983 2188 33992
rect 2136 33949 2145 33983
rect 2145 33949 2179 33983
rect 2179 33949 2188 33983
rect 2136 33940 2188 33949
rect 3240 33940 3292 33992
rect 3976 33940 4028 33992
rect 4620 33872 4672 33924
rect 2320 33847 2372 33856
rect 2320 33813 2329 33847
rect 2329 33813 2363 33847
rect 2363 33813 2372 33847
rect 2320 33804 2372 33813
rect 3056 33804 3108 33856
rect 4213 33702 4265 33754
rect 4277 33702 4329 33754
rect 4341 33702 4393 33754
rect 4405 33702 4457 33754
rect 4469 33702 4521 33754
rect 7477 33702 7529 33754
rect 7541 33702 7593 33754
rect 7605 33702 7657 33754
rect 7669 33702 7721 33754
rect 7733 33702 7785 33754
rect 3516 33600 3568 33652
rect 1584 33464 1636 33516
rect 2044 33464 2096 33516
rect 3424 33464 3476 33516
rect 9772 33464 9824 33516
rect 2136 33328 2188 33380
rect 3332 33328 3384 33380
rect 10048 33371 10100 33380
rect 10048 33337 10057 33371
rect 10057 33337 10091 33371
rect 10091 33337 10100 33371
rect 10048 33328 10100 33337
rect 1492 33260 1544 33312
rect 2320 33303 2372 33312
rect 2320 33269 2329 33303
rect 2329 33269 2363 33303
rect 2363 33269 2372 33303
rect 2320 33260 2372 33269
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5845 33158 5897 33210
rect 5909 33158 5961 33210
rect 5973 33158 6025 33210
rect 6037 33158 6089 33210
rect 6101 33158 6153 33210
rect 9109 33158 9161 33210
rect 9173 33158 9225 33210
rect 9237 33158 9289 33210
rect 9301 33158 9353 33210
rect 9365 33158 9417 33210
rect 9864 33056 9916 33108
rect 9680 32988 9732 33040
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 1952 32852 2004 32904
rect 2964 32852 3016 32904
rect 3240 32852 3292 32904
rect 3700 32852 3752 32904
rect 4068 32784 4120 32836
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 1676 32716 1728 32768
rect 1952 32716 2004 32768
rect 2320 32759 2372 32768
rect 2320 32725 2329 32759
rect 2329 32725 2363 32759
rect 2363 32725 2372 32759
rect 2320 32716 2372 32725
rect 3700 32716 3752 32768
rect 3884 32716 3936 32768
rect 10048 32759 10100 32768
rect 10048 32725 10057 32759
rect 10057 32725 10091 32759
rect 10091 32725 10100 32759
rect 10048 32716 10100 32725
rect 4213 32614 4265 32666
rect 4277 32614 4329 32666
rect 4341 32614 4393 32666
rect 4405 32614 4457 32666
rect 4469 32614 4521 32666
rect 7477 32614 7529 32666
rect 7541 32614 7593 32666
rect 7605 32614 7657 32666
rect 7669 32614 7721 32666
rect 7733 32614 7785 32666
rect 9772 32512 9824 32564
rect 3976 32444 4028 32496
rect 2044 32376 2096 32428
rect 2412 32376 2464 32428
rect 3240 32376 3292 32428
rect 1768 32308 1820 32360
rect 1492 32215 1544 32224
rect 1492 32181 1501 32215
rect 1501 32181 1535 32215
rect 1535 32181 1544 32215
rect 1492 32172 1544 32181
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5845 32070 5897 32122
rect 5909 32070 5961 32122
rect 5973 32070 6025 32122
rect 6037 32070 6089 32122
rect 6101 32070 6153 32122
rect 9109 32070 9161 32122
rect 9173 32070 9225 32122
rect 9237 32070 9289 32122
rect 9301 32070 9353 32122
rect 9365 32070 9417 32122
rect 5264 31968 5316 32020
rect 2780 31900 2832 31952
rect 10048 31943 10100 31952
rect 10048 31909 10057 31943
rect 10057 31909 10091 31943
rect 10091 31909 10100 31943
rect 10048 31900 10100 31909
rect 3792 31832 3844 31884
rect 2504 31807 2556 31816
rect 2504 31773 2513 31807
rect 2513 31773 2547 31807
rect 2547 31773 2556 31807
rect 2504 31764 2556 31773
rect 2504 31628 2556 31680
rect 3148 31628 3200 31680
rect 4213 31526 4265 31578
rect 4277 31526 4329 31578
rect 4341 31526 4393 31578
rect 4405 31526 4457 31578
rect 4469 31526 4521 31578
rect 7477 31526 7529 31578
rect 7541 31526 7593 31578
rect 7605 31526 7657 31578
rect 7669 31526 7721 31578
rect 7733 31526 7785 31578
rect 6644 31424 6696 31476
rect 296 31356 348 31408
rect 3056 31288 3108 31340
rect 3424 31220 3476 31272
rect 2136 31084 2188 31136
rect 2412 31084 2464 31136
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5845 30982 5897 31034
rect 5909 30982 5961 31034
rect 5973 30982 6025 31034
rect 6037 30982 6089 31034
rect 6101 30982 6153 31034
rect 9109 30982 9161 31034
rect 9173 30982 9225 31034
rect 9237 30982 9289 31034
rect 9301 30982 9353 31034
rect 9365 30982 9417 31034
rect 388 30880 440 30932
rect 3516 30880 3568 30932
rect 3792 30923 3844 30932
rect 3792 30889 3801 30923
rect 3801 30889 3835 30923
rect 3835 30889 3844 30923
rect 3792 30880 3844 30889
rect 1676 30812 1728 30864
rect 8668 30812 8720 30864
rect 2596 30744 2648 30796
rect 7104 30744 7156 30796
rect 3516 30676 3568 30728
rect 3976 30719 4028 30728
rect 3976 30685 3985 30719
rect 3985 30685 4019 30719
rect 4019 30685 4028 30719
rect 3976 30676 4028 30685
rect 9496 30676 9548 30728
rect 2964 30608 3016 30660
rect 10048 30583 10100 30592
rect 10048 30549 10057 30583
rect 10057 30549 10091 30583
rect 10091 30549 10100 30583
rect 10048 30540 10100 30549
rect 4213 30438 4265 30490
rect 4277 30438 4329 30490
rect 4341 30438 4393 30490
rect 4405 30438 4457 30490
rect 4469 30438 4521 30490
rect 7477 30438 7529 30490
rect 7541 30438 7593 30490
rect 7605 30438 7657 30490
rect 7669 30438 7721 30490
rect 7733 30438 7785 30490
rect 3148 30336 3200 30388
rect 2596 30268 2648 30320
rect 1676 30243 1728 30252
rect 1676 30209 1685 30243
rect 1685 30209 1719 30243
rect 1719 30209 1728 30243
rect 1676 30200 1728 30209
rect 2228 30243 2280 30252
rect 2228 30209 2237 30243
rect 2237 30209 2271 30243
rect 2271 30209 2280 30243
rect 2228 30200 2280 30209
rect 5356 30268 5408 30320
rect 2136 30132 2188 30184
rect 1492 30107 1544 30116
rect 1492 30073 1501 30107
rect 1501 30073 1535 30107
rect 1535 30073 1544 30107
rect 1492 30064 1544 30073
rect 3884 30064 3936 30116
rect 3056 29996 3108 30048
rect 10140 30039 10192 30048
rect 10140 30005 10149 30039
rect 10149 30005 10183 30039
rect 10183 30005 10192 30039
rect 10140 29996 10192 30005
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5845 29894 5897 29946
rect 5909 29894 5961 29946
rect 5973 29894 6025 29946
rect 6037 29894 6089 29946
rect 6101 29894 6153 29946
rect 9109 29894 9161 29946
rect 9173 29894 9225 29946
rect 9237 29894 9289 29946
rect 9301 29894 9353 29946
rect 9365 29894 9417 29946
rect 112 29792 164 29844
rect 3424 29792 3476 29844
rect 2136 29724 2188 29776
rect 1308 29656 1360 29708
rect 1584 29631 1636 29640
rect 1584 29597 1593 29631
rect 1593 29597 1627 29631
rect 1627 29597 1636 29631
rect 1584 29588 1636 29597
rect 480 29520 532 29572
rect 1768 29520 1820 29572
rect 3240 29631 3292 29640
rect 3240 29597 3249 29631
rect 3249 29597 3283 29631
rect 3283 29597 3292 29631
rect 3240 29588 3292 29597
rect 3424 29588 3476 29640
rect 3976 29631 4028 29640
rect 3976 29597 3985 29631
rect 3985 29597 4019 29631
rect 4019 29597 4028 29631
rect 3976 29588 4028 29597
rect 4712 29520 4764 29572
rect 3884 29452 3936 29504
rect 4620 29452 4672 29504
rect 4213 29350 4265 29402
rect 4277 29350 4329 29402
rect 4341 29350 4393 29402
rect 4405 29350 4457 29402
rect 4469 29350 4521 29402
rect 7477 29350 7529 29402
rect 7541 29350 7593 29402
rect 7605 29350 7657 29402
rect 7669 29350 7721 29402
rect 7733 29350 7785 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 1308 29180 1360 29232
rect 2964 29248 3016 29300
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 1584 29112 1636 29164
rect 2136 29112 2188 29164
rect 5080 29180 5132 29232
rect 3240 29155 3292 29164
rect 1768 29044 1820 29096
rect 3240 29121 3249 29155
rect 3249 29121 3283 29155
rect 3283 29121 3292 29155
rect 3240 29112 3292 29121
rect 2136 28976 2188 29028
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5845 28806 5897 28858
rect 5909 28806 5961 28858
rect 5973 28806 6025 28858
rect 6037 28806 6089 28858
rect 6101 28806 6153 28858
rect 9109 28806 9161 28858
rect 9173 28806 9225 28858
rect 9237 28806 9289 28858
rect 9301 28806 9353 28858
rect 9365 28806 9417 28858
rect 2320 28747 2372 28756
rect 2320 28713 2329 28747
rect 2329 28713 2363 28747
rect 2363 28713 2372 28747
rect 2320 28704 2372 28713
rect 3056 28747 3108 28756
rect 3056 28713 3065 28747
rect 3065 28713 3099 28747
rect 3099 28713 3108 28747
rect 3056 28704 3108 28713
rect 2504 28636 2556 28688
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 2872 28543 2924 28552
rect 2872 28509 2881 28543
rect 2881 28509 2915 28543
rect 2915 28509 2924 28543
rect 2872 28500 2924 28509
rect 3240 28432 3292 28484
rect 10140 28407 10192 28416
rect 10140 28373 10149 28407
rect 10149 28373 10183 28407
rect 10183 28373 10192 28407
rect 10140 28364 10192 28373
rect 4213 28262 4265 28314
rect 4277 28262 4329 28314
rect 4341 28262 4393 28314
rect 4405 28262 4457 28314
rect 4469 28262 4521 28314
rect 7477 28262 7529 28314
rect 7541 28262 7593 28314
rect 7605 28262 7657 28314
rect 7669 28262 7721 28314
rect 7733 28262 7785 28314
rect 1676 28160 1728 28212
rect 1768 28160 1820 28212
rect 2412 28067 2464 28076
rect 2412 28033 2421 28067
rect 2421 28033 2455 28067
rect 2455 28033 2464 28067
rect 2412 28024 2464 28033
rect 2964 27956 3016 28008
rect 1676 27888 1728 27940
rect 2044 27888 2096 27940
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5845 27718 5897 27770
rect 5909 27718 5961 27770
rect 5973 27718 6025 27770
rect 6037 27718 6089 27770
rect 6101 27718 6153 27770
rect 9109 27718 9161 27770
rect 9173 27718 9225 27770
rect 9237 27718 9289 27770
rect 9301 27718 9353 27770
rect 9365 27718 9417 27770
rect 940 27548 992 27600
rect 2964 27548 3016 27600
rect 3424 27480 3476 27532
rect 3976 27480 4028 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 2964 27455 3016 27464
rect 2964 27421 2973 27455
rect 2973 27421 3007 27455
rect 3007 27421 3016 27455
rect 2964 27412 3016 27421
rect 4620 27412 4672 27464
rect 5172 27412 5224 27464
rect 2136 27276 2188 27328
rect 2504 27276 2556 27328
rect 10140 27319 10192 27328
rect 10140 27285 10149 27319
rect 10149 27285 10183 27319
rect 10183 27285 10192 27319
rect 10140 27276 10192 27285
rect 4213 27174 4265 27226
rect 4277 27174 4329 27226
rect 4341 27174 4393 27226
rect 4405 27174 4457 27226
rect 4469 27174 4521 27226
rect 7477 27174 7529 27226
rect 7541 27174 7593 27226
rect 7605 27174 7657 27226
rect 7669 27174 7721 27226
rect 7733 27174 7785 27226
rect 848 27004 900 27056
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 3148 26979 3200 26988
rect 3148 26945 3157 26979
rect 3157 26945 3191 26979
rect 3191 26945 3200 26979
rect 3148 26936 3200 26945
rect 1860 26800 1912 26852
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5845 26630 5897 26682
rect 5909 26630 5961 26682
rect 5973 26630 6025 26682
rect 6037 26630 6089 26682
rect 6101 26630 6153 26682
rect 9109 26630 9161 26682
rect 9173 26630 9225 26682
rect 9237 26630 9289 26682
rect 9301 26630 9353 26682
rect 9365 26630 9417 26682
rect 1492 26571 1544 26580
rect 1492 26537 1501 26571
rect 1501 26537 1535 26571
rect 1535 26537 1544 26571
rect 1492 26528 1544 26537
rect 2504 26528 2556 26580
rect 572 26460 624 26512
rect 2688 26392 2740 26444
rect 10140 26435 10192 26444
rect 10140 26401 10149 26435
rect 10149 26401 10183 26435
rect 10183 26401 10192 26435
rect 10140 26392 10192 26401
rect 1768 26324 1820 26376
rect 2228 26367 2280 26376
rect 2228 26333 2237 26367
rect 2237 26333 2271 26367
rect 2271 26333 2280 26367
rect 2228 26324 2280 26333
rect 3056 26367 3108 26376
rect 3056 26333 3065 26367
rect 3065 26333 3099 26367
rect 3099 26333 3108 26367
rect 3056 26324 3108 26333
rect 3332 26256 3384 26308
rect 4213 26086 4265 26138
rect 4277 26086 4329 26138
rect 4341 26086 4393 26138
rect 4405 26086 4457 26138
rect 4469 26086 4521 26138
rect 7477 26086 7529 26138
rect 7541 26086 7593 26138
rect 7605 26086 7657 26138
rect 7669 26086 7721 26138
rect 7733 26086 7785 26138
rect 2228 26027 2280 26036
rect 2228 25993 2237 26027
rect 2237 25993 2271 26027
rect 2271 25993 2280 26027
rect 2228 25984 2280 25993
rect 2688 26027 2740 26036
rect 2688 25993 2697 26027
rect 2697 25993 2731 26027
rect 2731 25993 2740 26027
rect 2688 25984 2740 25993
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 1492 25848 1544 25900
rect 2872 25891 2924 25900
rect 2872 25857 2881 25891
rect 2881 25857 2915 25891
rect 2915 25857 2924 25891
rect 2872 25848 2924 25857
rect 2136 25644 2188 25696
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5845 25542 5897 25594
rect 5909 25542 5961 25594
rect 5973 25542 6025 25594
rect 6037 25542 6089 25594
rect 6101 25542 6153 25594
rect 9109 25542 9161 25594
rect 9173 25542 9225 25594
rect 9237 25542 9289 25594
rect 9301 25542 9353 25594
rect 9365 25542 9417 25594
rect 3700 25440 3752 25492
rect 10140 25483 10192 25492
rect 10140 25449 10149 25483
rect 10149 25449 10183 25483
rect 10183 25449 10192 25483
rect 10140 25440 10192 25449
rect 2780 25236 2832 25288
rect 4213 24998 4265 25050
rect 4277 24998 4329 25050
rect 4341 24998 4393 25050
rect 4405 24998 4457 25050
rect 4469 24998 4521 25050
rect 7477 24998 7529 25050
rect 7541 24998 7593 25050
rect 7605 24998 7657 25050
rect 7669 24998 7721 25050
rect 7733 24998 7785 25050
rect 1492 24760 1544 24812
rect 2136 24803 2188 24812
rect 2136 24769 2145 24803
rect 2145 24769 2179 24803
rect 2179 24769 2188 24803
rect 2136 24760 2188 24769
rect 2964 24803 3016 24812
rect 2964 24769 2973 24803
rect 2973 24769 3007 24803
rect 3007 24769 3016 24803
rect 2964 24760 3016 24769
rect 10140 24803 10192 24812
rect 10140 24769 10149 24803
rect 10149 24769 10183 24803
rect 10183 24769 10192 24803
rect 10140 24760 10192 24769
rect 1952 24692 2004 24744
rect 3240 24624 3292 24676
rect 3424 24556 3476 24608
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5845 24454 5897 24506
rect 5909 24454 5961 24506
rect 5973 24454 6025 24506
rect 6037 24454 6089 24506
rect 6101 24454 6153 24506
rect 9109 24454 9161 24506
rect 9173 24454 9225 24506
rect 9237 24454 9289 24506
rect 9301 24454 9353 24506
rect 9365 24454 9417 24506
rect 1216 24352 1268 24404
rect 3976 24284 4028 24336
rect 1676 24216 1728 24268
rect 3424 24216 3476 24268
rect 3976 24191 4028 24200
rect 3976 24157 3985 24191
rect 3985 24157 4019 24191
rect 4019 24157 4028 24191
rect 3976 24148 4028 24157
rect 2320 24080 2372 24132
rect 2504 24080 2556 24132
rect 3240 24012 3292 24064
rect 3700 24012 3752 24064
rect 4213 23910 4265 23962
rect 4277 23910 4329 23962
rect 4341 23910 4393 23962
rect 4405 23910 4457 23962
rect 4469 23910 4521 23962
rect 7477 23910 7529 23962
rect 7541 23910 7593 23962
rect 7605 23910 7657 23962
rect 7669 23910 7721 23962
rect 7733 23910 7785 23962
rect 1216 23672 1268 23724
rect 1952 23672 2004 23724
rect 2412 23740 2464 23792
rect 2504 23672 2556 23724
rect 3240 23715 3292 23724
rect 3240 23681 3249 23715
rect 3249 23681 3283 23715
rect 3283 23681 3292 23715
rect 3240 23672 3292 23681
rect 9864 23715 9916 23724
rect 3424 23604 3476 23656
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 1400 23468 1452 23520
rect 7380 23536 7432 23588
rect 8944 23468 8996 23520
rect 10048 23511 10100 23520
rect 10048 23477 10057 23511
rect 10057 23477 10091 23511
rect 10091 23477 10100 23511
rect 10048 23468 10100 23477
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5845 23366 5897 23418
rect 5909 23366 5961 23418
rect 5973 23366 6025 23418
rect 6037 23366 6089 23418
rect 6101 23366 6153 23418
rect 9109 23366 9161 23418
rect 9173 23366 9225 23418
rect 9237 23366 9289 23418
rect 9301 23366 9353 23418
rect 9365 23366 9417 23418
rect 3884 23264 3936 23316
rect 9864 23264 9916 23316
rect 10140 23307 10192 23316
rect 10140 23273 10149 23307
rect 10149 23273 10183 23307
rect 10183 23273 10192 23307
rect 10140 23264 10192 23273
rect 2872 23196 2924 23248
rect 3424 23196 3476 23248
rect 2688 23128 2740 23180
rect 1676 23103 1728 23112
rect 1676 23069 1685 23103
rect 1685 23069 1719 23103
rect 1719 23069 1728 23103
rect 1676 23060 1728 23069
rect 2412 23060 2464 23112
rect 2964 23060 3016 23112
rect 3240 22992 3292 23044
rect 4620 22924 4672 22976
rect 4213 22822 4265 22874
rect 4277 22822 4329 22874
rect 4341 22822 4393 22874
rect 4405 22822 4457 22874
rect 4469 22822 4521 22874
rect 7477 22822 7529 22874
rect 7541 22822 7593 22874
rect 7605 22822 7657 22874
rect 7669 22822 7721 22874
rect 7733 22822 7785 22874
rect 2228 22720 2280 22772
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 2136 22584 2188 22636
rect 2504 22720 2556 22772
rect 3056 22720 3108 22772
rect 3424 22720 3476 22772
rect 3516 22720 3568 22772
rect 2872 22652 2924 22704
rect 6276 22652 6328 22704
rect 3424 22584 3476 22636
rect 9772 22584 9824 22636
rect 2504 22516 2556 22568
rect 2412 22448 2464 22500
rect 2688 22448 2740 22500
rect 10048 22491 10100 22500
rect 10048 22457 10057 22491
rect 10057 22457 10091 22491
rect 10091 22457 10100 22491
rect 10048 22448 10100 22457
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5845 22278 5897 22330
rect 5909 22278 5961 22330
rect 5973 22278 6025 22330
rect 6037 22278 6089 22330
rect 6101 22278 6153 22330
rect 9109 22278 9161 22330
rect 9173 22278 9225 22330
rect 9237 22278 9289 22330
rect 9301 22278 9353 22330
rect 9365 22278 9417 22330
rect 3056 22176 3108 22228
rect 3792 22176 3844 22228
rect 1124 22040 1176 22092
rect 2320 22015 2372 22024
rect 2320 21981 2329 22015
rect 2329 21981 2363 22015
rect 2363 21981 2372 22015
rect 2320 21972 2372 21981
rect 2412 22015 2464 22024
rect 2412 21981 2421 22015
rect 2421 21981 2455 22015
rect 2455 21981 2464 22015
rect 3148 22015 3200 22024
rect 2412 21972 2464 21981
rect 3148 21981 3157 22015
rect 3157 21981 3191 22015
rect 3191 21981 3200 22015
rect 3148 21972 3200 21981
rect 4804 21904 4856 21956
rect 9864 22015 9916 22024
rect 9864 21981 9873 22015
rect 9873 21981 9907 22015
rect 9907 21981 9916 22015
rect 9864 21972 9916 21981
rect 7288 21836 7340 21888
rect 9772 21836 9824 21888
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 4213 21734 4265 21786
rect 4277 21734 4329 21786
rect 4341 21734 4393 21786
rect 4405 21734 4457 21786
rect 4469 21734 4521 21786
rect 7477 21734 7529 21786
rect 7541 21734 7593 21786
rect 7605 21734 7657 21786
rect 7669 21734 7721 21786
rect 7733 21734 7785 21786
rect 2964 21675 3016 21684
rect 2964 21641 2973 21675
rect 2973 21641 3007 21675
rect 3007 21641 3016 21675
rect 2964 21632 3016 21641
rect 1492 21564 1544 21616
rect 4804 21564 4856 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 3056 21496 3108 21548
rect 9772 21496 9824 21548
rect 2228 21360 2280 21412
rect 2504 21292 2556 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5845 21190 5897 21242
rect 5909 21190 5961 21242
rect 5973 21190 6025 21242
rect 6037 21190 6089 21242
rect 6101 21190 6153 21242
rect 9109 21190 9161 21242
rect 9173 21190 9225 21242
rect 9237 21190 9289 21242
rect 9301 21190 9353 21242
rect 9365 21190 9417 21242
rect 1032 21088 1084 21140
rect 3700 21088 3752 21140
rect 4068 21088 4120 21140
rect 9864 21131 9916 21140
rect 9864 21097 9873 21131
rect 9873 21097 9907 21131
rect 9907 21097 9916 21131
rect 9864 21088 9916 21097
rect 2504 20884 2556 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 3148 20816 3200 20868
rect 3792 20816 3844 20868
rect 4068 20748 4120 20800
rect 4213 20646 4265 20698
rect 4277 20646 4329 20698
rect 4341 20646 4393 20698
rect 4405 20646 4457 20698
rect 4469 20646 4521 20698
rect 7477 20646 7529 20698
rect 7541 20646 7593 20698
rect 7605 20646 7657 20698
rect 7669 20646 7721 20698
rect 7733 20646 7785 20698
rect 3148 20587 3200 20596
rect 3148 20553 3157 20587
rect 3157 20553 3191 20587
rect 3191 20553 3200 20587
rect 3148 20544 3200 20553
rect 2780 20408 2832 20460
rect 9680 20408 9732 20460
rect 2964 20340 3016 20392
rect 3424 20272 3476 20324
rect 10048 20315 10100 20324
rect 10048 20281 10057 20315
rect 10057 20281 10091 20315
rect 10091 20281 10100 20315
rect 10048 20272 10100 20281
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5845 20102 5897 20154
rect 5909 20102 5961 20154
rect 5973 20102 6025 20154
rect 6037 20102 6089 20154
rect 6101 20102 6153 20154
rect 9109 20102 9161 20154
rect 9173 20102 9225 20154
rect 9237 20102 9289 20154
rect 9301 20102 9353 20154
rect 9365 20102 9417 20154
rect 3792 20000 3844 20052
rect 2780 19796 2832 19848
rect 3148 19839 3200 19848
rect 3148 19805 3157 19839
rect 3157 19805 3191 19839
rect 3191 19805 3200 19839
rect 3148 19796 3200 19805
rect 9864 19839 9916 19848
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 1860 19660 1912 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 4213 19558 4265 19610
rect 4277 19558 4329 19610
rect 4341 19558 4393 19610
rect 4405 19558 4457 19610
rect 4469 19558 4521 19610
rect 7477 19558 7529 19610
rect 7541 19558 7593 19610
rect 7605 19558 7657 19610
rect 7669 19558 7721 19610
rect 7733 19558 7785 19610
rect 9772 19456 9824 19508
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 2964 19320 3016 19372
rect 3608 19184 3660 19236
rect 2504 19159 2556 19168
rect 2504 19125 2513 19159
rect 2513 19125 2547 19159
rect 2547 19125 2556 19159
rect 2504 19116 2556 19125
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5845 19014 5897 19066
rect 5909 19014 5961 19066
rect 5973 19014 6025 19066
rect 6037 19014 6089 19066
rect 6101 19014 6153 19066
rect 9109 19014 9161 19066
rect 9173 19014 9225 19066
rect 9237 19014 9289 19066
rect 9301 19014 9353 19066
rect 9365 19014 9417 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 9864 18912 9916 18964
rect 2136 18776 2188 18828
rect 4068 18776 4120 18828
rect 2412 18751 2464 18760
rect 2412 18717 2421 18751
rect 2421 18717 2455 18751
rect 2455 18717 2464 18751
rect 2412 18708 2464 18717
rect 2688 18708 2740 18760
rect 3976 18751 4028 18760
rect 3976 18717 3985 18751
rect 3985 18717 4019 18751
rect 4019 18717 4028 18751
rect 3976 18708 4028 18717
rect 9772 18708 9824 18760
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 4213 18470 4265 18522
rect 4277 18470 4329 18522
rect 4341 18470 4393 18522
rect 4405 18470 4457 18522
rect 4469 18470 4521 18522
rect 7477 18470 7529 18522
rect 7541 18470 7593 18522
rect 7605 18470 7657 18522
rect 7669 18470 7721 18522
rect 7733 18470 7785 18522
rect 1676 18411 1728 18420
rect 1676 18377 1685 18411
rect 1685 18377 1719 18411
rect 1719 18377 1728 18411
rect 1676 18368 1728 18377
rect 2412 18411 2464 18420
rect 2412 18377 2421 18411
rect 2421 18377 2455 18411
rect 2455 18377 2464 18411
rect 2412 18368 2464 18377
rect 9680 18368 9732 18420
rect 2228 18300 2280 18352
rect 3056 18300 3108 18352
rect 2412 18232 2464 18284
rect 2688 18232 2740 18284
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 3792 18164 3844 18216
rect 1860 18096 1912 18148
rect 9956 18232 10008 18284
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5845 17926 5897 17978
rect 5909 17926 5961 17978
rect 5973 17926 6025 17978
rect 6037 17926 6089 17978
rect 6101 17926 6153 17978
rect 9109 17926 9161 17978
rect 9173 17926 9225 17978
rect 9237 17926 9289 17978
rect 9301 17926 9353 17978
rect 9365 17926 9417 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 3792 17867 3844 17876
rect 3792 17833 3801 17867
rect 3801 17833 3835 17867
rect 3835 17833 3844 17867
rect 3792 17824 3844 17833
rect 1584 17756 1636 17808
rect 3240 17688 3292 17740
rect 2504 17663 2556 17672
rect 2504 17629 2513 17663
rect 2513 17629 2547 17663
rect 2547 17629 2556 17663
rect 2504 17620 2556 17629
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 9864 17663 9916 17672
rect 9864 17629 9873 17663
rect 9873 17629 9907 17663
rect 9907 17629 9916 17663
rect 9864 17620 9916 17629
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 4213 17382 4265 17434
rect 4277 17382 4329 17434
rect 4341 17382 4393 17434
rect 4405 17382 4457 17434
rect 4469 17382 4521 17434
rect 7477 17382 7529 17434
rect 7541 17382 7593 17434
rect 7605 17382 7657 17434
rect 7669 17382 7721 17434
rect 7733 17382 7785 17434
rect 9956 17323 10008 17332
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 1492 17144 1544 17196
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 1768 16940 1820 16992
rect 2228 16940 2280 16992
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5845 16838 5897 16890
rect 5909 16838 5961 16890
rect 5973 16838 6025 16890
rect 6037 16838 6089 16890
rect 6101 16838 6153 16890
rect 9109 16838 9161 16890
rect 9173 16838 9225 16890
rect 9237 16838 9289 16890
rect 9301 16838 9353 16890
rect 9365 16838 9417 16890
rect 2228 16600 2280 16652
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 2320 16464 2372 16516
rect 2504 16464 2556 16516
rect 9680 16532 9732 16584
rect 2596 16439 2648 16448
rect 2596 16405 2605 16439
rect 2605 16405 2639 16439
rect 2639 16405 2648 16439
rect 2596 16396 2648 16405
rect 9772 16396 9824 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 4213 16294 4265 16346
rect 4277 16294 4329 16346
rect 4341 16294 4393 16346
rect 4405 16294 4457 16346
rect 4469 16294 4521 16346
rect 7477 16294 7529 16346
rect 7541 16294 7593 16346
rect 7605 16294 7657 16346
rect 7669 16294 7721 16346
rect 7733 16294 7785 16346
rect 2136 16192 2188 16244
rect 1676 16124 1728 16176
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 2320 16056 2372 16108
rect 2044 15988 2096 16040
rect 3240 15988 3292 16040
rect 1676 15852 1728 15904
rect 2596 15920 2648 15972
rect 2412 15852 2464 15904
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5845 15750 5897 15802
rect 5909 15750 5961 15802
rect 5973 15750 6025 15802
rect 6037 15750 6089 15802
rect 6101 15750 6153 15802
rect 9109 15750 9161 15802
rect 9173 15750 9225 15802
rect 9237 15750 9289 15802
rect 9301 15750 9353 15802
rect 9365 15750 9417 15802
rect 1676 15648 1728 15700
rect 2044 15648 2096 15700
rect 9864 15648 9916 15700
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 2504 15376 2556 15428
rect 1584 15308 1636 15360
rect 1768 15308 1820 15360
rect 4213 15206 4265 15258
rect 4277 15206 4329 15258
rect 4341 15206 4393 15258
rect 4405 15206 4457 15258
rect 4469 15206 4521 15258
rect 7477 15206 7529 15258
rect 7541 15206 7593 15258
rect 7605 15206 7657 15258
rect 7669 15206 7721 15258
rect 7733 15206 7785 15258
rect 1400 15104 1452 15156
rect 2136 15104 2188 15156
rect 3056 15104 3108 15156
rect 1584 15036 1636 15088
rect 1860 14968 1912 15020
rect 2136 14832 2188 14884
rect 2964 14968 3016 15020
rect 2412 14900 2464 14952
rect 10048 14875 10100 14884
rect 10048 14841 10057 14875
rect 10057 14841 10091 14875
rect 10091 14841 10100 14875
rect 10048 14832 10100 14841
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5845 14662 5897 14714
rect 5909 14662 5961 14714
rect 5973 14662 6025 14714
rect 6037 14662 6089 14714
rect 6101 14662 6153 14714
rect 9109 14662 9161 14714
rect 9173 14662 9225 14714
rect 9237 14662 9289 14714
rect 9301 14662 9353 14714
rect 9365 14662 9417 14714
rect 1492 14560 1544 14612
rect 1676 14492 1728 14544
rect 1492 14424 1544 14476
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 1676 14356 1728 14408
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 4213 14118 4265 14170
rect 4277 14118 4329 14170
rect 4341 14118 4393 14170
rect 4405 14118 4457 14170
rect 4469 14118 4521 14170
rect 7477 14118 7529 14170
rect 7541 14118 7593 14170
rect 7605 14118 7657 14170
rect 7669 14118 7721 14170
rect 7733 14118 7785 14170
rect 1492 14016 1544 14068
rect 2964 14016 3016 14068
rect 9680 14016 9732 14068
rect 2320 13948 2372 14000
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 3148 13812 3200 13864
rect 10140 13812 10192 13864
rect 10048 13719 10100 13728
rect 10048 13685 10057 13719
rect 10057 13685 10091 13719
rect 10091 13685 10100 13719
rect 10048 13676 10100 13685
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5845 13574 5897 13626
rect 5909 13574 5961 13626
rect 5973 13574 6025 13626
rect 6037 13574 6089 13626
rect 6101 13574 6153 13626
rect 9109 13574 9161 13626
rect 9173 13574 9225 13626
rect 9237 13574 9289 13626
rect 9301 13574 9353 13626
rect 9365 13574 9417 13626
rect 3240 13404 3292 13456
rect 2044 13336 2096 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 1768 13200 1820 13252
rect 2044 13200 2096 13252
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 4213 13030 4265 13082
rect 4277 13030 4329 13082
rect 4341 13030 4393 13082
rect 4405 13030 4457 13082
rect 4469 13030 4521 13082
rect 7477 13030 7529 13082
rect 7541 13030 7593 13082
rect 7605 13030 7657 13082
rect 7669 13030 7721 13082
rect 7733 13030 7785 13082
rect 1492 12928 1544 12980
rect 1768 12928 1820 12980
rect 7840 12928 7892 12980
rect 2228 12792 2280 12844
rect 3424 12792 3476 12844
rect 9772 12792 9824 12844
rect 1308 12724 1360 12776
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5845 12486 5897 12538
rect 5909 12486 5961 12538
rect 5973 12486 6025 12538
rect 6037 12486 6089 12538
rect 6101 12486 6153 12538
rect 9109 12486 9161 12538
rect 9173 12486 9225 12538
rect 9237 12486 9289 12538
rect 9301 12486 9353 12538
rect 9365 12486 9417 12538
rect 7932 12384 7984 12436
rect 2044 12248 2096 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 3884 12112 3936 12164
rect 9772 12044 9824 12096
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 4213 11942 4265 11994
rect 4277 11942 4329 11994
rect 4341 11942 4393 11994
rect 4405 11942 4457 11994
rect 4469 11942 4521 11994
rect 7477 11942 7529 11994
rect 7541 11942 7593 11994
rect 7605 11942 7657 11994
rect 7669 11942 7721 11994
rect 7733 11942 7785 11994
rect 7196 11840 7248 11892
rect 3240 11772 3292 11824
rect 1768 11704 1820 11756
rect 2228 11704 2280 11756
rect 3424 11747 3476 11756
rect 3424 11713 3433 11747
rect 3433 11713 3467 11747
rect 3467 11713 3476 11747
rect 3424 11704 3476 11713
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 1308 11636 1360 11688
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 9864 11500 9916 11552
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5845 11398 5897 11450
rect 5909 11398 5961 11450
rect 5973 11398 6025 11450
rect 6037 11398 6089 11450
rect 6101 11398 6153 11450
rect 9109 11398 9161 11450
rect 9173 11398 9225 11450
rect 9237 11398 9289 11450
rect 9301 11398 9353 11450
rect 9365 11398 9417 11450
rect 3608 11296 3660 11348
rect 9680 11228 9732 11280
rect 1492 11160 1544 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2228 11092 2280 11144
rect 3884 11092 3936 11144
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 9772 11024 9824 11076
rect 4213 10854 4265 10906
rect 4277 10854 4329 10906
rect 4341 10854 4393 10906
rect 4405 10854 4457 10906
rect 4469 10854 4521 10906
rect 7477 10854 7529 10906
rect 7541 10854 7593 10906
rect 7605 10854 7657 10906
rect 7669 10854 7721 10906
rect 7733 10854 7785 10906
rect 9036 10684 9088 10736
rect 2136 10616 2188 10668
rect 3056 10616 3108 10668
rect 1308 10548 1360 10600
rect 2964 10480 3016 10532
rect 3976 10616 4028 10668
rect 9680 10616 9732 10668
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5845 10310 5897 10362
rect 5909 10310 5961 10362
rect 5973 10310 6025 10362
rect 6037 10310 6089 10362
rect 6101 10310 6153 10362
rect 9109 10310 9161 10362
rect 9173 10310 9225 10362
rect 9237 10310 9289 10362
rect 9301 10310 9353 10362
rect 9365 10310 9417 10362
rect 3148 10072 3200 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2136 10004 2188 10056
rect 4620 10004 4672 10056
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 9864 9868 9916 9920
rect 4213 9766 4265 9818
rect 4277 9766 4329 9818
rect 4341 9766 4393 9818
rect 4405 9766 4457 9818
rect 4469 9766 4521 9818
rect 7477 9766 7529 9818
rect 7541 9766 7593 9818
rect 7605 9766 7657 9818
rect 7669 9766 7721 9818
rect 7733 9766 7785 9818
rect 3976 9664 4028 9716
rect 10140 9664 10192 9716
rect 3700 9596 3752 9648
rect 2320 9528 2372 9580
rect 2412 9528 2464 9580
rect 3240 9528 3292 9580
rect 4620 9528 4672 9580
rect 9772 9528 9824 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2504 9392 2556 9444
rect 10048 9435 10100 9444
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5845 9222 5897 9274
rect 5909 9222 5961 9274
rect 5973 9222 6025 9274
rect 6037 9222 6089 9274
rect 6101 9222 6153 9274
rect 9109 9222 9161 9274
rect 9173 9222 9225 9274
rect 9237 9222 9289 9274
rect 9301 9222 9353 9274
rect 9365 9222 9417 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 6552 9052 6604 9104
rect 2412 8984 2464 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2872 8916 2924 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3148 8916 3200 8968
rect 3516 8916 3568 8968
rect 9864 8959 9916 8968
rect 9864 8925 9873 8959
rect 9873 8925 9907 8959
rect 9907 8925 9916 8959
rect 9864 8916 9916 8925
rect 1584 8848 1636 8900
rect 6460 8848 6512 8900
rect 6184 8780 6236 8832
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 4213 8678 4265 8730
rect 4277 8678 4329 8730
rect 4341 8678 4393 8730
rect 4405 8678 4457 8730
rect 4469 8678 4521 8730
rect 7477 8678 7529 8730
rect 7541 8678 7593 8730
rect 7605 8678 7657 8730
rect 7669 8678 7721 8730
rect 7733 8678 7785 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 6736 8508 6788 8560
rect 1492 8440 1544 8492
rect 1584 8440 1636 8492
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 3700 8372 3752 8424
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5845 8134 5897 8186
rect 5909 8134 5961 8186
rect 5973 8134 6025 8186
rect 6037 8134 6089 8186
rect 6101 8134 6153 8186
rect 9109 8134 9161 8186
rect 9173 8134 9225 8186
rect 9237 8134 9289 8186
rect 9301 8134 9353 8186
rect 9365 8134 9417 8186
rect 3976 8075 4028 8084
rect 3976 8041 3985 8075
rect 3985 8041 4019 8075
rect 4019 8041 4028 8075
rect 3976 8032 4028 8041
rect 2780 7964 2832 8016
rect 3792 7964 3844 8016
rect 2412 7896 2464 7948
rect 3148 7896 3200 7948
rect 3424 7896 3476 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 1860 7828 1912 7880
rect 2504 7828 2556 7880
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 9864 7760 9916 7812
rect 4213 7590 4265 7642
rect 4277 7590 4329 7642
rect 4341 7590 4393 7642
rect 4405 7590 4457 7642
rect 4469 7590 4521 7642
rect 7477 7590 7529 7642
rect 7541 7590 7593 7642
rect 7605 7590 7657 7642
rect 7669 7590 7721 7642
rect 7733 7590 7785 7642
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 1216 7420 1268 7472
rect 2044 7352 2096 7404
rect 3608 7352 3660 7404
rect 9864 7395 9916 7404
rect 9864 7361 9873 7395
rect 9873 7361 9907 7395
rect 9907 7361 9916 7395
rect 9864 7352 9916 7361
rect 3700 7284 3752 7336
rect 9864 7148 9916 7200
rect 10048 7191 10100 7200
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5845 7046 5897 7098
rect 5909 7046 5961 7098
rect 5973 7046 6025 7098
rect 6037 7046 6089 7098
rect 6101 7046 6153 7098
rect 9109 7046 9161 7098
rect 9173 7046 9225 7098
rect 9237 7046 9289 7098
rect 9301 7046 9353 7098
rect 9365 7046 9417 7098
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1492 6740 1544 6792
rect 4068 6672 4120 6724
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 4213 6502 4265 6554
rect 4277 6502 4329 6554
rect 4341 6502 4393 6554
rect 4405 6502 4457 6554
rect 4469 6502 4521 6554
rect 7477 6502 7529 6554
rect 7541 6502 7593 6554
rect 7605 6502 7657 6554
rect 7669 6502 7721 6554
rect 7733 6502 7785 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 3516 6443 3568 6452
rect 3516 6409 3525 6443
rect 3525 6409 3559 6443
rect 3559 6409 3568 6443
rect 3516 6400 3568 6409
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2964 6264 3016 6316
rect 3332 6307 3384 6316
rect 3332 6273 3341 6307
rect 3341 6273 3375 6307
rect 3375 6273 3384 6307
rect 3332 6264 3384 6273
rect 3884 6128 3936 6180
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5845 5958 5897 6010
rect 5909 5958 5961 6010
rect 5973 5958 6025 6010
rect 6037 5958 6089 6010
rect 6101 5958 6153 6010
rect 9109 5958 9161 6010
rect 9173 5958 9225 6010
rect 9237 5958 9289 6010
rect 9301 5958 9353 6010
rect 9365 5958 9417 6010
rect 1492 5856 1544 5908
rect 1308 5652 1360 5704
rect 1584 5652 1636 5704
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 4213 5414 4265 5466
rect 4277 5414 4329 5466
rect 4341 5414 4393 5466
rect 4405 5414 4457 5466
rect 4469 5414 4521 5466
rect 7477 5414 7529 5466
rect 7541 5414 7593 5466
rect 7605 5414 7657 5466
rect 7669 5414 7721 5466
rect 7733 5414 7785 5466
rect 5540 5312 5592 5364
rect 1584 5176 1636 5228
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 3240 5244 3292 5296
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 3608 5219 3660 5228
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 4712 5108 4764 5160
rect 2964 5015 3016 5024
rect 2964 4981 2973 5015
rect 2973 4981 3007 5015
rect 3007 4981 3016 5015
rect 2964 4972 3016 4981
rect 4160 4972 4212 5024
rect 7104 4972 7156 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5845 4870 5897 4922
rect 5909 4870 5961 4922
rect 5973 4870 6025 4922
rect 6037 4870 6089 4922
rect 6101 4870 6153 4922
rect 9109 4870 9161 4922
rect 9173 4870 9225 4922
rect 9237 4870 9289 4922
rect 9301 4870 9353 4922
rect 9365 4870 9417 4922
rect 3424 4768 3476 4820
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 4160 4768 4212 4820
rect 9864 4768 9916 4820
rect 4712 4700 4764 4752
rect 2964 4632 3016 4684
rect 9772 4632 9824 4684
rect 3424 4564 3476 4616
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 7104 4564 7156 4616
rect 3792 4496 3844 4548
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 4213 4326 4265 4378
rect 4277 4326 4329 4378
rect 4341 4326 4393 4378
rect 4405 4326 4457 4378
rect 4469 4326 4521 4378
rect 7477 4326 7529 4378
rect 7541 4326 7593 4378
rect 7605 4326 7657 4378
rect 7669 4326 7721 4378
rect 7733 4326 7785 4378
rect 1952 4156 2004 4208
rect 3608 4156 3660 4208
rect 3516 4088 3568 4140
rect 3148 3952 3200 4004
rect 4620 4020 4672 4072
rect 5540 3952 5592 4004
rect 8024 3884 8076 3936
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5845 3782 5897 3834
rect 5909 3782 5961 3834
rect 5973 3782 6025 3834
rect 6037 3782 6089 3834
rect 6101 3782 6153 3834
rect 9109 3782 9161 3834
rect 9173 3782 9225 3834
rect 9237 3782 9289 3834
rect 9301 3782 9353 3834
rect 9365 3782 9417 3834
rect 2504 3680 2556 3732
rect 3148 3544 3200 3596
rect 2228 3476 2280 3528
rect 3516 3476 3568 3528
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 7932 3408 7984 3460
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 4213 3238 4265 3290
rect 4277 3238 4329 3290
rect 4341 3238 4393 3290
rect 4405 3238 4457 3290
rect 4469 3238 4521 3290
rect 7477 3238 7529 3290
rect 7541 3238 7593 3290
rect 7605 3238 7657 3290
rect 7669 3238 7721 3290
rect 7733 3238 7785 3290
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 3424 3179 3476 3188
rect 3424 3145 3433 3179
rect 3433 3145 3467 3179
rect 3467 3145 3476 3179
rect 3424 3136 3476 3145
rect 3700 3136 3752 3188
rect 2412 3000 2464 3052
rect 3608 3043 3660 3052
rect 3608 3009 3617 3043
rect 3617 3009 3651 3043
rect 3651 3009 3660 3043
rect 3608 3000 3660 3009
rect 4160 3000 4212 3052
rect 8024 3000 8076 3052
rect 9772 3000 9824 3052
rect 5080 2932 5132 2984
rect 9864 2864 9916 2916
rect 5632 2796 5684 2848
rect 9496 2796 9548 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5845 2694 5897 2746
rect 5909 2694 5961 2746
rect 5973 2694 6025 2746
rect 6037 2694 6089 2746
rect 6101 2694 6153 2746
rect 9109 2694 9161 2746
rect 9173 2694 9225 2746
rect 9237 2694 9289 2746
rect 9301 2694 9353 2746
rect 9365 2694 9417 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2320 2592 2372 2644
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4620 2592 4672 2644
rect 5080 2635 5132 2644
rect 5080 2601 5089 2635
rect 5089 2601 5123 2635
rect 5123 2601 5132 2635
rect 5080 2592 5132 2601
rect 2412 2524 2464 2576
rect 1400 2431 1452 2440
rect 1400 2397 1409 2431
rect 1409 2397 1443 2431
rect 1443 2397 1452 2431
rect 1400 2388 1452 2397
rect 2780 2388 2832 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 3976 2431 4028 2440
rect 2872 2388 2924 2397
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5540 2388 5592 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 4213 2150 4265 2202
rect 4277 2150 4329 2202
rect 4341 2150 4393 2202
rect 4405 2150 4457 2202
rect 4469 2150 4521 2202
rect 7477 2150 7529 2202
rect 7541 2150 7593 2202
rect 7605 2150 7657 2202
rect 7669 2150 7721 2202
rect 7733 2150 7785 2202
rect 2872 1028 2924 1080
rect 5264 1028 5316 1080
rect 2780 484 2832 536
rect 4620 484 4672 536
<< metal2 >>
rect 2962 79656 3018 79665
rect 2962 79591 3018 79600
rect 1398 79248 1454 79257
rect 1398 79183 1454 79192
rect 1412 77586 1440 79183
rect 2778 78840 2834 78849
rect 2778 78775 2834 78784
rect 2792 78130 2820 78775
rect 2780 78124 2832 78130
rect 2780 78066 2832 78072
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 1400 77580 1452 77586
rect 1400 77522 1452 77528
rect 2976 77518 3004 79591
rect 10046 79520 10102 79529
rect 10046 79455 10102 79464
rect 3514 78432 3570 78441
rect 3514 78367 3570 78376
rect 3422 77616 3478 77625
rect 3422 77551 3478 77560
rect 2964 77512 3016 77518
rect 2964 77454 3016 77460
rect 2136 77376 2188 77382
rect 2136 77318 2188 77324
rect 1400 77036 1452 77042
rect 1400 76978 1452 76984
rect 112 76560 164 76566
rect 112 76502 164 76508
rect 124 60734 152 76502
rect 1412 76430 1440 76978
rect 1400 76424 1452 76430
rect 1400 76366 1452 76372
rect 1952 76424 2004 76430
rect 1952 76366 2004 76372
rect 1768 76084 1820 76090
rect 1768 76026 1820 76032
rect 1492 75948 1544 75954
rect 1492 75890 1544 75896
rect 1400 74860 1452 74866
rect 1400 74802 1452 74808
rect 1412 74361 1440 74802
rect 1504 74497 1532 75890
rect 1676 74860 1728 74866
rect 1676 74802 1728 74808
rect 1584 74656 1636 74662
rect 1584 74598 1636 74604
rect 1490 74488 1546 74497
rect 1490 74423 1546 74432
rect 1398 74352 1454 74361
rect 1398 74287 1454 74296
rect 1400 74248 1452 74254
rect 1400 74190 1452 74196
rect 572 73568 624 73574
rect 572 73510 624 73516
rect 388 67244 440 67250
rect 388 67186 440 67192
rect 204 61804 256 61810
rect 204 61746 256 61752
rect 32 60706 152 60734
rect 32 48346 60 60706
rect 112 57588 164 57594
rect 112 57530 164 57536
rect 20 48340 72 48346
rect 20 48282 72 48288
rect 124 46186 152 57530
rect 32 46158 152 46186
rect 32 39506 60 46158
rect 112 46096 164 46102
rect 112 46038 164 46044
rect 20 39500 72 39506
rect 20 39442 72 39448
rect 124 29850 152 46038
rect 216 41682 244 61746
rect 296 52964 348 52970
rect 296 52906 348 52912
rect 204 41676 256 41682
rect 204 41618 256 41624
rect 204 41540 256 41546
rect 204 41482 256 41488
rect 216 36582 244 41482
rect 204 36576 256 36582
rect 204 36518 256 36524
rect 308 31414 336 52906
rect 400 49162 428 67186
rect 480 60512 532 60518
rect 480 60454 532 60460
rect 492 54806 520 60454
rect 480 54800 532 54806
rect 480 54742 532 54748
rect 480 51808 532 51814
rect 480 51750 532 51756
rect 388 49156 440 49162
rect 388 49098 440 49104
rect 388 48884 440 48890
rect 388 48826 440 48832
rect 400 46306 428 48826
rect 388 46300 440 46306
rect 388 46242 440 46248
rect 492 46186 520 51750
rect 400 46158 520 46186
rect 296 31408 348 31414
rect 296 31350 348 31356
rect 400 30938 428 46158
rect 480 46096 532 46102
rect 480 46038 532 46044
rect 388 30932 440 30938
rect 388 30874 440 30880
rect 112 29844 164 29850
rect 112 29786 164 29792
rect 492 29578 520 46038
rect 584 43994 612 73510
rect 1412 73273 1440 74190
rect 1492 74112 1544 74118
rect 1492 74054 1544 74060
rect 1398 73264 1454 73273
rect 1398 73199 1454 73208
rect 1504 72842 1532 74054
rect 1136 72814 1532 72842
rect 1136 69442 1164 72814
rect 1400 72684 1452 72690
rect 1400 72626 1452 72632
rect 1216 72072 1268 72078
rect 1216 72014 1268 72020
rect 1228 71097 1256 72014
rect 1412 71913 1440 72626
rect 1492 71936 1544 71942
rect 1398 71904 1454 71913
rect 1492 71878 1544 71884
rect 1398 71839 1454 71848
rect 1308 71596 1360 71602
rect 1308 71538 1360 71544
rect 1214 71088 1270 71097
rect 1214 71023 1270 71032
rect 1216 70916 1268 70922
rect 1216 70858 1268 70864
rect 1228 70496 1256 70858
rect 1320 70689 1348 71538
rect 1400 70984 1452 70990
rect 1400 70926 1452 70932
rect 1306 70680 1362 70689
rect 1306 70615 1362 70624
rect 1308 70508 1360 70514
rect 1228 70468 1308 70496
rect 1308 70450 1360 70456
rect 1320 69884 1348 70450
rect 1412 70281 1440 70926
rect 1398 70272 1454 70281
rect 1398 70207 1454 70216
rect 1400 69896 1452 69902
rect 1320 69856 1400 69884
rect 1400 69838 1452 69844
rect 1412 69562 1440 69838
rect 1400 69556 1452 69562
rect 1400 69498 1452 69504
rect 1136 69414 1440 69442
rect 1308 69352 1360 69358
rect 1308 69294 1360 69300
rect 1216 69216 1268 69222
rect 1216 69158 1268 69164
rect 1032 68332 1084 68338
rect 1032 68274 1084 68280
rect 940 63368 992 63374
rect 940 63310 992 63316
rect 848 62280 900 62286
rect 848 62222 900 62228
rect 664 58676 716 58682
rect 664 58618 716 58624
rect 572 43988 624 43994
rect 572 43930 624 43936
rect 572 43716 624 43722
rect 572 43658 624 43664
rect 584 43178 612 43658
rect 572 43172 624 43178
rect 572 43114 624 43120
rect 584 36718 612 43114
rect 676 40730 704 58618
rect 756 56840 808 56846
rect 756 56782 808 56788
rect 664 40724 716 40730
rect 664 40666 716 40672
rect 768 38010 796 56782
rect 860 42566 888 62222
rect 952 43382 980 63310
rect 1044 50250 1072 68274
rect 1124 67788 1176 67794
rect 1124 67730 1176 67736
rect 1032 50244 1084 50250
rect 1032 50186 1084 50192
rect 1136 49774 1164 67730
rect 1228 60518 1256 69158
rect 1320 68785 1348 69294
rect 1412 69018 1440 69414
rect 1400 69012 1452 69018
rect 1400 68954 1452 68960
rect 1400 68808 1452 68814
rect 1306 68776 1362 68785
rect 1400 68750 1452 68756
rect 1306 68711 1362 68720
rect 1308 68264 1360 68270
rect 1308 68206 1360 68212
rect 1320 67697 1348 68206
rect 1412 68105 1440 68750
rect 1398 68096 1454 68105
rect 1398 68031 1454 68040
rect 1400 67720 1452 67726
rect 1306 67688 1362 67697
rect 1400 67662 1452 67668
rect 1306 67623 1362 67632
rect 1412 67289 1440 67662
rect 1398 67280 1454 67289
rect 1398 67215 1454 67224
rect 1400 67176 1452 67182
rect 1400 67118 1452 67124
rect 1412 66881 1440 67118
rect 1398 66872 1454 66881
rect 1398 66807 1454 66816
rect 1400 66632 1452 66638
rect 1400 66574 1452 66580
rect 1412 66337 1440 66574
rect 1398 66328 1454 66337
rect 1308 66292 1360 66298
rect 1398 66263 1454 66272
rect 1308 66234 1360 66240
rect 1320 64410 1348 66234
rect 1398 65920 1454 65929
rect 1398 65855 1454 65864
rect 1412 65550 1440 65855
rect 1504 65600 1532 71878
rect 1596 69902 1624 74598
rect 1688 73778 1716 74802
rect 1676 73772 1728 73778
rect 1676 73714 1728 73720
rect 1688 73166 1716 73714
rect 1676 73160 1728 73166
rect 1676 73102 1728 73108
rect 1688 72690 1716 73102
rect 1676 72684 1728 72690
rect 1676 72626 1728 72632
rect 1676 72480 1728 72486
rect 1676 72422 1728 72428
rect 1584 69896 1636 69902
rect 1584 69838 1636 69844
rect 1584 69760 1636 69766
rect 1584 69702 1636 69708
rect 1596 68474 1624 69702
rect 1584 68468 1636 68474
rect 1584 68410 1636 68416
rect 1688 68354 1716 72422
rect 1780 70650 1808 76026
rect 1964 75954 1992 76366
rect 1952 75948 2004 75954
rect 1952 75890 2004 75896
rect 1964 75342 1992 75890
rect 1952 75336 2004 75342
rect 1952 75278 2004 75284
rect 1964 73778 1992 75278
rect 1952 73772 2004 73778
rect 1952 73714 2004 73720
rect 1952 73568 2004 73574
rect 1952 73510 2004 73516
rect 1860 73092 1912 73098
rect 1860 73034 1912 73040
rect 1872 72826 1900 73034
rect 1860 72820 1912 72826
rect 1860 72762 1912 72768
rect 1860 71392 1912 71398
rect 1860 71334 1912 71340
rect 1768 70644 1820 70650
rect 1768 70586 1820 70592
rect 1768 70508 1820 70514
rect 1768 70450 1820 70456
rect 1780 69902 1808 70450
rect 1768 69896 1820 69902
rect 1768 69838 1820 69844
rect 1780 69426 1808 69838
rect 1768 69420 1820 69426
rect 1768 69362 1820 69368
rect 1780 68882 1808 69362
rect 1768 68876 1820 68882
rect 1768 68818 1820 68824
rect 1768 68672 1820 68678
rect 1768 68614 1820 68620
rect 1596 68326 1716 68354
rect 1596 66230 1624 68326
rect 1676 68196 1728 68202
rect 1676 68138 1728 68144
rect 1688 66298 1716 68138
rect 1780 66473 1808 68614
rect 1872 67634 1900 71334
rect 1964 69494 1992 73510
rect 2042 72448 2098 72457
rect 2042 72383 2098 72392
rect 2056 72078 2084 72383
rect 2044 72072 2096 72078
rect 2044 72014 2096 72020
rect 2044 71732 2096 71738
rect 2044 71674 2096 71680
rect 2056 71058 2084 71674
rect 2044 71052 2096 71058
rect 2044 70994 2096 71000
rect 2044 70848 2096 70854
rect 2044 70790 2096 70796
rect 1952 69488 2004 69494
rect 1952 69430 2004 69436
rect 1952 69012 2004 69018
rect 1952 68954 2004 68960
rect 1964 68406 1992 68954
rect 1952 68400 2004 68406
rect 1952 68342 2004 68348
rect 1872 67606 1992 67634
rect 1860 66632 1912 66638
rect 1860 66574 1912 66580
rect 1766 66464 1822 66473
rect 1766 66399 1822 66408
rect 1676 66292 1728 66298
rect 1676 66234 1728 66240
rect 1584 66224 1636 66230
rect 1584 66166 1636 66172
rect 1674 66192 1730 66201
rect 1674 66127 1676 66136
rect 1728 66127 1730 66136
rect 1676 66098 1728 66104
rect 1768 65680 1820 65686
rect 1766 65648 1768 65657
rect 1820 65648 1822 65657
rect 1676 65612 1728 65618
rect 1504 65572 1624 65600
rect 1400 65544 1452 65550
rect 1400 65486 1452 65492
rect 1492 64456 1544 64462
rect 1320 64404 1492 64410
rect 1320 64398 1544 64404
rect 1320 64382 1532 64398
rect 1400 63776 1452 63782
rect 1400 63718 1452 63724
rect 1412 62529 1440 63718
rect 1492 63232 1544 63238
rect 1492 63174 1544 63180
rect 1398 62520 1454 62529
rect 1398 62455 1454 62464
rect 1400 62348 1452 62354
rect 1400 62290 1452 62296
rect 1412 62234 1440 62290
rect 1320 62206 1440 62234
rect 1216 60512 1268 60518
rect 1216 60454 1268 60460
rect 1216 60240 1268 60246
rect 1216 60182 1268 60188
rect 1228 55418 1256 60182
rect 1320 58970 1348 62206
rect 1400 62144 1452 62150
rect 1504 62121 1532 63174
rect 1596 62966 1624 65572
rect 1766 65583 1822 65592
rect 1676 65554 1728 65560
rect 1584 62960 1636 62966
rect 1584 62902 1636 62908
rect 1400 62086 1452 62092
rect 1490 62112 1546 62121
rect 1412 61169 1440 62086
rect 1490 62047 1546 62056
rect 1492 61736 1544 61742
rect 1490 61704 1492 61713
rect 1544 61704 1546 61713
rect 1490 61639 1546 61648
rect 1492 61600 1544 61606
rect 1492 61542 1544 61548
rect 1398 61160 1454 61169
rect 1398 61095 1454 61104
rect 1400 61056 1452 61062
rect 1400 60998 1452 61004
rect 1412 59945 1440 60998
rect 1504 60761 1532 61542
rect 1688 60790 1716 65554
rect 1768 65408 1820 65414
rect 1768 65350 1820 65356
rect 1676 60784 1728 60790
rect 1490 60752 1546 60761
rect 1676 60726 1728 60732
rect 1490 60687 1546 60696
rect 1676 60648 1728 60654
rect 1676 60590 1728 60596
rect 1688 60110 1716 60590
rect 1676 60104 1728 60110
rect 1676 60046 1728 60052
rect 1398 59936 1454 59945
rect 1398 59871 1454 59880
rect 1688 59770 1716 60046
rect 1676 59764 1728 59770
rect 1676 59706 1728 59712
rect 1492 59424 1544 59430
rect 1492 59366 1544 59372
rect 1400 59220 1452 59226
rect 1400 59162 1452 59168
rect 1412 59129 1440 59162
rect 1398 59120 1454 59129
rect 1398 59055 1454 59064
rect 1320 58942 1440 58970
rect 1308 58880 1360 58886
rect 1308 58822 1360 58828
rect 1320 58478 1348 58822
rect 1308 58472 1360 58478
rect 1308 58414 1360 58420
rect 1320 58002 1348 58414
rect 1308 57996 1360 58002
rect 1308 57938 1360 57944
rect 1412 56506 1440 58942
rect 1504 58585 1532 59366
rect 1584 59152 1636 59158
rect 1584 59094 1636 59100
rect 1596 59022 1624 59094
rect 1688 59090 1716 59706
rect 1676 59084 1728 59090
rect 1676 59026 1728 59032
rect 1584 59016 1636 59022
rect 1584 58958 1636 58964
rect 1582 58848 1638 58857
rect 1582 58783 1638 58792
rect 1490 58576 1546 58585
rect 1490 58511 1546 58520
rect 1492 57248 1544 57254
rect 1492 57190 1544 57196
rect 1504 56953 1532 57190
rect 1490 56944 1546 56953
rect 1490 56879 1546 56888
rect 1492 56704 1544 56710
rect 1492 56646 1544 56652
rect 1504 56545 1532 56646
rect 1490 56536 1546 56545
rect 1400 56500 1452 56506
rect 1490 56471 1546 56480
rect 1400 56442 1452 56448
rect 1400 56296 1452 56302
rect 1320 56244 1400 56250
rect 1320 56238 1452 56244
rect 1320 56222 1440 56238
rect 1216 55412 1268 55418
rect 1216 55354 1268 55360
rect 1320 55162 1348 56222
rect 1400 56160 1452 56166
rect 1400 56102 1452 56108
rect 1412 55321 1440 56102
rect 1492 55616 1544 55622
rect 1492 55558 1544 55564
rect 1504 55457 1532 55558
rect 1490 55448 1546 55457
rect 1490 55383 1546 55392
rect 1596 55350 1624 58783
rect 1674 58576 1730 58585
rect 1674 58511 1676 58520
rect 1728 58511 1730 58520
rect 1676 58482 1728 58488
rect 1688 58002 1716 58482
rect 1676 57996 1728 58002
rect 1676 57938 1728 57944
rect 1676 56500 1728 56506
rect 1676 56442 1728 56448
rect 1584 55344 1636 55350
rect 1398 55312 1454 55321
rect 1584 55286 1636 55292
rect 1398 55247 1454 55256
rect 1584 55208 1636 55214
rect 1320 55156 1584 55162
rect 1320 55150 1636 55156
rect 1320 55134 1624 55150
rect 1216 54868 1268 54874
rect 1216 54810 1268 54816
rect 1124 49768 1176 49774
rect 1124 49710 1176 49716
rect 1032 47116 1084 47122
rect 1032 47058 1084 47064
rect 940 43376 992 43382
rect 940 43318 992 43324
rect 940 43240 992 43246
rect 940 43182 992 43188
rect 848 42560 900 42566
rect 848 42502 900 42508
rect 952 42378 980 43182
rect 860 42350 980 42378
rect 756 38004 808 38010
rect 756 37946 808 37952
rect 572 36712 624 36718
rect 572 36654 624 36660
rect 572 36576 624 36582
rect 572 36518 624 36524
rect 480 29572 532 29578
rect 480 29514 532 29520
rect 584 26518 612 36518
rect 756 36236 808 36242
rect 756 36178 808 36184
rect 572 26512 624 26518
rect 572 26454 624 26460
rect 768 26234 796 36178
rect 860 27062 888 42350
rect 1044 41414 1072 47058
rect 1124 46708 1176 46714
rect 1124 46650 1176 46656
rect 1136 43246 1164 46650
rect 1228 46102 1256 54810
rect 1400 54528 1452 54534
rect 1400 54470 1452 54476
rect 1412 53961 1440 54470
rect 1492 53984 1544 53990
rect 1398 53952 1454 53961
rect 1492 53926 1544 53932
rect 1398 53887 1454 53896
rect 1308 53576 1360 53582
rect 1504 53553 1532 53926
rect 1596 53786 1624 55134
rect 1584 53780 1636 53786
rect 1584 53722 1636 53728
rect 1308 53518 1360 53524
rect 1490 53544 1546 53553
rect 1320 52018 1348 53518
rect 1490 53479 1546 53488
rect 1400 52896 1452 52902
rect 1400 52838 1452 52844
rect 1412 52193 1440 52838
rect 1492 52352 1544 52358
rect 1492 52294 1544 52300
rect 1398 52184 1454 52193
rect 1398 52119 1454 52128
rect 1308 52012 1360 52018
rect 1308 51954 1360 51960
rect 1320 50522 1348 51954
rect 1504 51785 1532 52294
rect 1596 51882 1624 53722
rect 1688 52034 1716 56442
rect 1780 53718 1808 65350
rect 1768 53712 1820 53718
rect 1768 53654 1820 53660
rect 1872 53564 1900 66574
rect 1964 65618 1992 67606
rect 1952 65612 2004 65618
rect 1952 65554 2004 65560
rect 2056 65498 2084 70790
rect 2148 69306 2176 77318
rect 3436 77042 3464 77551
rect 2228 77036 2280 77042
rect 2228 76978 2280 76984
rect 2964 77036 3016 77042
rect 2964 76978 3016 76984
rect 3332 77036 3384 77042
rect 3332 76978 3384 76984
rect 3424 77036 3476 77042
rect 3424 76978 3476 76984
rect 2240 76430 2268 76978
rect 2412 76832 2464 76838
rect 2412 76774 2464 76780
rect 2228 76424 2280 76430
rect 2228 76366 2280 76372
rect 2240 75886 2268 76366
rect 2228 75880 2280 75886
rect 2228 75822 2280 75828
rect 2240 75342 2268 75822
rect 2228 75336 2280 75342
rect 2228 75278 2280 75284
rect 2240 74866 2268 75278
rect 2228 74860 2280 74866
rect 2228 74802 2280 74808
rect 2228 73772 2280 73778
rect 2228 73714 2280 73720
rect 2240 73234 2268 73714
rect 2228 73228 2280 73234
rect 2228 73170 2280 73176
rect 2228 73024 2280 73030
rect 2228 72966 2280 72972
rect 2240 72554 2268 72966
rect 2320 72684 2372 72690
rect 2320 72626 2372 72632
rect 2228 72548 2280 72554
rect 2228 72490 2280 72496
rect 2332 72434 2360 72626
rect 2240 72406 2360 72434
rect 2240 71738 2268 72406
rect 2320 71936 2372 71942
rect 2320 71878 2372 71884
rect 2228 71732 2280 71738
rect 2228 71674 2280 71680
rect 2228 71596 2280 71602
rect 2228 71538 2280 71544
rect 2240 71505 2268 71538
rect 2226 71496 2282 71505
rect 2226 71431 2282 71440
rect 2228 71392 2280 71398
rect 2228 71334 2280 71340
rect 2240 69766 2268 71334
rect 2228 69760 2280 69766
rect 2228 69702 2280 69708
rect 2148 69278 2268 69306
rect 2136 69216 2188 69222
rect 2136 69158 2188 69164
rect 1964 65470 2084 65498
rect 1964 58546 1992 65470
rect 2044 65068 2096 65074
rect 2044 65010 2096 65016
rect 2056 64462 2084 65010
rect 2148 64977 2176 69158
rect 2240 66502 2268 69278
rect 2332 66570 2360 71878
rect 2424 70990 2452 76774
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 2976 76265 3004 76978
rect 3056 76832 3108 76838
rect 3056 76774 3108 76780
rect 3240 76832 3292 76838
rect 3240 76774 3292 76780
rect 2962 76256 3018 76265
rect 2962 76191 3018 76200
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2964 75200 3016 75206
rect 2964 75142 3016 75148
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2976 73846 3004 75142
rect 2964 73840 3016 73846
rect 2964 73782 3016 73788
rect 2780 73772 2832 73778
rect 2780 73714 2832 73720
rect 2792 73681 2820 73714
rect 2778 73672 2834 73681
rect 2778 73607 2834 73616
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2964 73228 3016 73234
rect 2964 73170 3016 73176
rect 2780 73160 2832 73166
rect 2780 73102 2832 73108
rect 2504 73024 2556 73030
rect 2504 72966 2556 72972
rect 2412 70984 2464 70990
rect 2412 70926 2464 70932
rect 2412 70644 2464 70650
rect 2412 70586 2464 70592
rect 2320 66564 2372 66570
rect 2320 66506 2372 66512
rect 2228 66496 2280 66502
rect 2228 66438 2280 66444
rect 2228 66088 2280 66094
rect 2228 66030 2280 66036
rect 2240 65074 2268 66030
rect 2228 65068 2280 65074
rect 2228 65010 2280 65016
rect 2134 64968 2190 64977
rect 2134 64903 2190 64912
rect 2136 64864 2188 64870
rect 2136 64806 2188 64812
rect 2044 64456 2096 64462
rect 2044 64398 2096 64404
rect 2056 63458 2084 64398
rect 2148 63594 2176 64806
rect 2228 64456 2280 64462
rect 2228 64398 2280 64404
rect 2240 64054 2268 64398
rect 2228 64048 2280 64054
rect 2228 63990 2280 63996
rect 2228 63776 2280 63782
rect 2226 63744 2228 63753
rect 2280 63744 2282 63753
rect 2226 63679 2282 63688
rect 2424 63594 2452 70586
rect 2516 66314 2544 72966
rect 2792 72865 2820 73102
rect 2778 72856 2834 72865
rect 2778 72791 2834 72800
rect 2976 72690 3004 73170
rect 2964 72684 3016 72690
rect 2964 72626 3016 72632
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2596 70984 2648 70990
rect 2596 70926 2648 70932
rect 2608 70514 2636 70926
rect 2976 70854 3004 72626
rect 3068 72622 3096 76774
rect 3148 76424 3200 76430
rect 3148 76366 3200 76372
rect 3160 75857 3188 76366
rect 3252 76090 3280 76774
rect 3344 76537 3372 76978
rect 3330 76528 3386 76537
rect 3330 76463 3386 76472
rect 3528 76430 3556 78367
rect 4620 78124 4672 78130
rect 4620 78066 4672 78072
rect 4066 78024 4122 78033
rect 4066 77959 4122 77968
rect 3608 77580 3660 77586
rect 3608 77522 3660 77528
rect 3516 76424 3568 76430
rect 3516 76366 3568 76372
rect 3424 76288 3476 76294
rect 3424 76230 3476 76236
rect 3240 76084 3292 76090
rect 3240 76026 3292 76032
rect 3332 76084 3384 76090
rect 3332 76026 3384 76032
rect 3146 75848 3202 75857
rect 3146 75783 3202 75792
rect 3240 75812 3292 75818
rect 3240 75754 3292 75760
rect 3148 75336 3200 75342
rect 3148 75278 3200 75284
rect 3160 75041 3188 75278
rect 3146 75032 3202 75041
rect 3146 74967 3202 74976
rect 3148 74860 3200 74866
rect 3148 74802 3200 74808
rect 3160 73234 3188 74802
rect 3148 73228 3200 73234
rect 3148 73170 3200 73176
rect 3056 72616 3108 72622
rect 3056 72558 3108 72564
rect 2964 70848 3016 70854
rect 2964 70790 3016 70796
rect 2596 70508 2648 70514
rect 2596 70450 2648 70456
rect 2964 70508 3016 70514
rect 2964 70450 3016 70456
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2976 69873 3004 70450
rect 3056 69896 3108 69902
rect 2962 69864 3018 69873
rect 3056 69838 3108 69844
rect 2962 69799 3018 69808
rect 2596 69760 2648 69766
rect 2596 69702 2648 69708
rect 2608 69290 2636 69702
rect 2964 69420 3016 69426
rect 2964 69362 3016 69368
rect 2596 69284 2648 69290
rect 2596 69226 2648 69232
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 2596 68944 2648 68950
rect 2596 68886 2648 68892
rect 2608 68270 2636 68886
rect 2872 68808 2924 68814
rect 2870 68776 2872 68785
rect 2924 68776 2926 68785
rect 2870 68711 2926 68720
rect 2780 68332 2832 68338
rect 2884 68320 2912 68711
rect 2976 68513 3004 69362
rect 3068 68921 3096 69838
rect 3054 68912 3110 68921
rect 3054 68847 3110 68856
rect 2962 68504 3018 68513
rect 2962 68439 3018 68448
rect 3056 68332 3108 68338
rect 2832 68292 3004 68320
rect 2780 68274 2832 68280
rect 2596 68264 2648 68270
rect 2596 68206 2648 68212
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2976 66756 3004 68292
rect 3056 68274 3108 68280
rect 2884 66728 3004 66756
rect 2516 66286 2636 66314
rect 2884 66298 2912 66728
rect 2964 66496 3016 66502
rect 2964 66438 3016 66444
rect 2608 66230 2636 66286
rect 2872 66292 2924 66298
rect 2872 66234 2924 66240
rect 2596 66224 2648 66230
rect 2596 66166 2648 66172
rect 2504 66156 2556 66162
rect 2504 66098 2556 66104
rect 2148 63566 2268 63594
rect 2056 63430 2176 63458
rect 2044 63368 2096 63374
rect 2044 63310 2096 63316
rect 2056 62354 2084 63310
rect 2148 62898 2176 63430
rect 2136 62892 2188 62898
rect 2136 62834 2188 62840
rect 2044 62348 2096 62354
rect 2044 62290 2096 62296
rect 2044 61804 2096 61810
rect 2044 61746 2096 61752
rect 1952 58540 2004 58546
rect 1952 58482 2004 58488
rect 1952 57928 2004 57934
rect 1952 57870 2004 57876
rect 1964 56302 1992 57870
rect 1952 56296 2004 56302
rect 1952 56238 2004 56244
rect 1952 56160 2004 56166
rect 1952 56102 2004 56108
rect 1964 53786 1992 56102
rect 2056 55944 2084 61746
rect 2148 60858 2176 62834
rect 2136 60852 2188 60858
rect 2136 60794 2188 60800
rect 2240 60734 2268 63566
rect 2148 60706 2268 60734
rect 2332 63566 2452 63594
rect 2516 65532 2544 66098
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2688 65544 2740 65550
rect 2516 65504 2688 65532
rect 2148 56166 2176 60706
rect 2228 60648 2280 60654
rect 2228 60590 2280 60596
rect 2240 57474 2268 60590
rect 2332 59702 2360 63566
rect 2516 63492 2544 65504
rect 2976 65521 3004 66438
rect 3068 66162 3096 68274
rect 3252 66774 3280 75754
rect 3344 72826 3372 76026
rect 3332 72820 3384 72826
rect 3332 72762 3384 72768
rect 3332 69420 3384 69426
rect 3332 69362 3384 69368
rect 3344 69329 3372 69362
rect 3330 69320 3386 69329
rect 3330 69255 3386 69264
rect 3436 68746 3464 76230
rect 3620 76106 3648 77522
rect 4080 77518 4108 77959
rect 3976 77512 4028 77518
rect 3976 77454 4028 77460
rect 4068 77512 4120 77518
rect 4068 77454 4120 77460
rect 3792 77376 3844 77382
rect 3792 77318 3844 77324
rect 3884 77376 3936 77382
rect 3884 77318 3936 77324
rect 3528 76078 3648 76106
rect 3528 75818 3556 76078
rect 3608 75948 3660 75954
rect 3608 75890 3660 75896
rect 3516 75812 3568 75818
rect 3516 75754 3568 75760
rect 3620 75449 3648 75890
rect 3606 75440 3662 75449
rect 3606 75375 3662 75384
rect 3804 74934 3832 77318
rect 3896 75410 3924 77318
rect 3988 77081 4016 77454
rect 4213 77276 4521 77296
rect 4213 77274 4219 77276
rect 4275 77274 4299 77276
rect 4355 77274 4379 77276
rect 4435 77274 4459 77276
rect 4515 77274 4521 77276
rect 4275 77222 4277 77274
rect 4457 77222 4459 77274
rect 4213 77220 4219 77222
rect 4275 77220 4299 77222
rect 4355 77220 4379 77222
rect 4435 77220 4459 77222
rect 4515 77220 4521 77222
rect 4213 77200 4521 77220
rect 3974 77072 4030 77081
rect 4632 77042 4660 78066
rect 9494 78024 9550 78033
rect 9494 77959 9550 77968
rect 5845 77820 6153 77840
rect 5845 77818 5851 77820
rect 5907 77818 5931 77820
rect 5987 77818 6011 77820
rect 6067 77818 6091 77820
rect 6147 77818 6153 77820
rect 5907 77766 5909 77818
rect 6089 77766 6091 77818
rect 5845 77764 5851 77766
rect 5907 77764 5931 77766
rect 5987 77764 6011 77766
rect 6067 77764 6091 77766
rect 6147 77764 6153 77766
rect 5845 77744 6153 77764
rect 9109 77820 9417 77840
rect 9109 77818 9115 77820
rect 9171 77818 9195 77820
rect 9251 77818 9275 77820
rect 9331 77818 9355 77820
rect 9411 77818 9417 77820
rect 9171 77766 9173 77818
rect 9353 77766 9355 77818
rect 9109 77764 9115 77766
rect 9171 77764 9195 77766
rect 9251 77764 9275 77766
rect 9331 77764 9355 77766
rect 9411 77764 9417 77766
rect 9109 77744 9417 77764
rect 9404 77512 9456 77518
rect 9404 77454 9456 77460
rect 5264 77376 5316 77382
rect 5264 77318 5316 77324
rect 3974 77007 4030 77016
rect 4620 77036 4672 77042
rect 4620 76978 4672 76984
rect 5276 76362 5304 77318
rect 7477 77276 7785 77296
rect 7477 77274 7483 77276
rect 7539 77274 7563 77276
rect 7619 77274 7643 77276
rect 7699 77274 7723 77276
rect 7779 77274 7785 77276
rect 7539 77222 7541 77274
rect 7721 77222 7723 77274
rect 7477 77220 7483 77222
rect 7539 77220 7563 77222
rect 7619 77220 7643 77222
rect 7699 77220 7723 77222
rect 7779 77220 7785 77222
rect 7477 77200 7785 77220
rect 9416 77217 9444 77454
rect 9402 77208 9458 77217
rect 9402 77143 9458 77152
rect 9508 77042 9536 77959
rect 10060 77518 10088 79455
rect 10966 78704 11022 78713
rect 10966 78639 10968 78648
rect 11020 78639 11022 78648
rect 10968 78610 11020 78616
rect 10048 77512 10100 77518
rect 10048 77454 10100 77460
rect 9496 77036 9548 77042
rect 9496 76978 9548 76984
rect 5540 76900 5592 76906
rect 5540 76842 5592 76848
rect 5264 76356 5316 76362
rect 5264 76298 5316 76304
rect 4213 76188 4521 76208
rect 4213 76186 4219 76188
rect 4275 76186 4299 76188
rect 4355 76186 4379 76188
rect 4435 76186 4459 76188
rect 4515 76186 4521 76188
rect 4275 76134 4277 76186
rect 4457 76134 4459 76186
rect 4213 76132 4219 76134
rect 4275 76132 4299 76134
rect 4355 76132 4379 76134
rect 4435 76132 4459 76134
rect 4515 76132 4521 76134
rect 4213 76112 4521 76132
rect 3976 75744 4028 75750
rect 3976 75686 4028 75692
rect 3884 75404 3936 75410
rect 3884 75346 3936 75352
rect 3792 74928 3844 74934
rect 3792 74870 3844 74876
rect 3608 70032 3660 70038
rect 3608 69974 3660 69980
rect 3516 69216 3568 69222
rect 3516 69158 3568 69164
rect 3424 68740 3476 68746
rect 3424 68682 3476 68688
rect 3240 66768 3292 66774
rect 3240 66710 3292 66716
rect 3240 66632 3292 66638
rect 3240 66574 3292 66580
rect 3148 66564 3200 66570
rect 3148 66506 3200 66512
rect 3056 66156 3108 66162
rect 3056 66098 3108 66104
rect 2688 65486 2740 65492
rect 2962 65512 3018 65521
rect 3068 65482 3096 66098
rect 3160 65686 3188 66506
rect 3148 65680 3200 65686
rect 3148 65622 3200 65628
rect 2962 65447 3018 65456
rect 3056 65476 3108 65482
rect 3056 65418 3108 65424
rect 3148 65476 3200 65482
rect 3148 65418 3200 65424
rect 3068 65074 3096 65418
rect 3056 65068 3108 65074
rect 3056 65010 3108 65016
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 2780 64320 2832 64326
rect 2778 64288 2780 64297
rect 2832 64288 2834 64297
rect 2778 64223 2834 64232
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2424 63464 2544 63492
rect 2872 63504 2924 63510
rect 2424 62354 2452 63464
rect 2872 63446 2924 63452
rect 2504 63368 2556 63374
rect 2504 63310 2556 63316
rect 2412 62348 2464 62354
rect 2412 62290 2464 62296
rect 2516 60897 2544 63310
rect 2884 62937 2912 63446
rect 3054 63336 3110 63345
rect 3054 63271 3110 63280
rect 3068 63238 3096 63271
rect 3056 63232 3108 63238
rect 3056 63174 3108 63180
rect 2870 62928 2926 62937
rect 2870 62863 2926 62872
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 2964 62280 3016 62286
rect 3160 62234 3188 65418
rect 2964 62222 3016 62228
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 2976 61334 3004 62222
rect 3068 62206 3188 62234
rect 2964 61328 3016 61334
rect 2964 61270 3016 61276
rect 2502 60888 2558 60897
rect 2502 60823 2558 60832
rect 2596 60852 2648 60858
rect 2596 60794 2648 60800
rect 2502 60752 2558 60761
rect 2502 60687 2558 60696
rect 2516 60602 2544 60687
rect 2424 60574 2544 60602
rect 2320 59696 2372 59702
rect 2320 59638 2372 59644
rect 2320 59560 2372 59566
rect 2320 59502 2372 59508
rect 2332 59022 2360 59502
rect 2320 59016 2372 59022
rect 2320 58958 2372 58964
rect 2332 58585 2360 58958
rect 2318 58576 2374 58585
rect 2318 58511 2374 58520
rect 2424 58426 2452 60574
rect 2608 60500 2636 60794
rect 3068 60734 3096 62206
rect 3148 61056 3200 61062
rect 3148 60998 3200 61004
rect 2976 60706 3096 60734
rect 2778 60616 2834 60625
rect 2778 60551 2780 60560
rect 2832 60551 2834 60560
rect 2780 60522 2832 60528
rect 2516 60472 2636 60500
rect 2516 60314 2544 60472
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2504 60308 2556 60314
rect 2504 60250 2556 60256
rect 2502 60208 2558 60217
rect 2502 60143 2558 60152
rect 2332 58398 2452 58426
rect 2332 57798 2360 58398
rect 2412 58336 2464 58342
rect 2412 58278 2464 58284
rect 2424 58177 2452 58278
rect 2410 58168 2466 58177
rect 2410 58103 2466 58112
rect 2412 58064 2464 58070
rect 2412 58006 2464 58012
rect 2320 57792 2372 57798
rect 2320 57734 2372 57740
rect 2240 57446 2360 57474
rect 2226 57352 2282 57361
rect 2226 57287 2228 57296
rect 2280 57287 2282 57296
rect 2228 57258 2280 57264
rect 2228 56704 2280 56710
rect 2228 56646 2280 56652
rect 2136 56160 2188 56166
rect 2136 56102 2188 56108
rect 2240 56001 2268 56646
rect 2226 55992 2282 56001
rect 2056 55916 2176 55944
rect 2226 55927 2282 55936
rect 2044 55072 2096 55078
rect 2044 55014 2096 55020
rect 1952 53780 2004 53786
rect 1952 53722 2004 53728
rect 1780 53536 1900 53564
rect 1780 52154 1808 53536
rect 1860 53440 1912 53446
rect 1860 53382 1912 53388
rect 1872 52578 1900 53382
rect 1952 53100 2004 53106
rect 1952 53042 2004 53048
rect 1964 52698 1992 53042
rect 1952 52692 2004 52698
rect 1952 52634 2004 52640
rect 1872 52550 1992 52578
rect 1860 52488 1912 52494
rect 1860 52430 1912 52436
rect 1768 52148 1820 52154
rect 1768 52090 1820 52096
rect 1688 52006 1808 52034
rect 1674 51912 1730 51921
rect 1584 51876 1636 51882
rect 1674 51847 1730 51856
rect 1584 51818 1636 51824
rect 1490 51776 1546 51785
rect 1490 51711 1546 51720
rect 1400 51264 1452 51270
rect 1400 51206 1452 51212
rect 1308 50516 1360 50522
rect 1308 50458 1360 50464
rect 1412 50425 1440 51206
rect 1492 50720 1544 50726
rect 1492 50662 1544 50668
rect 1398 50416 1454 50425
rect 1308 50380 1360 50386
rect 1398 50351 1454 50360
rect 1308 50322 1360 50328
rect 1320 48890 1348 50322
rect 1504 50017 1532 50662
rect 1596 50318 1624 51818
rect 1688 50454 1716 51847
rect 1676 50448 1728 50454
rect 1676 50390 1728 50396
rect 1584 50312 1636 50318
rect 1584 50254 1636 50260
rect 1490 50008 1546 50017
rect 1490 49943 1546 49952
rect 1596 49842 1624 50254
rect 1676 50176 1728 50182
rect 1676 50118 1728 50124
rect 1584 49836 1636 49842
rect 1584 49778 1636 49784
rect 1492 49700 1544 49706
rect 1492 49642 1544 49648
rect 1400 49632 1452 49638
rect 1400 49574 1452 49580
rect 1308 48884 1360 48890
rect 1308 48826 1360 48832
rect 1308 47660 1360 47666
rect 1308 47602 1360 47608
rect 1216 46096 1268 46102
rect 1216 46038 1268 46044
rect 1216 43988 1268 43994
rect 1216 43930 1268 43936
rect 1124 43240 1176 43246
rect 1124 43182 1176 43188
rect 1228 41478 1256 43930
rect 1216 41472 1268 41478
rect 1216 41414 1268 41420
rect 952 41386 1072 41414
rect 952 27606 980 41386
rect 1216 40928 1268 40934
rect 1216 40870 1268 40876
rect 1228 40225 1256 40870
rect 1214 40216 1270 40225
rect 1214 40151 1270 40160
rect 1216 39840 1268 39846
rect 1216 39782 1268 39788
rect 1228 38865 1256 39782
rect 1214 38856 1270 38865
rect 1214 38791 1270 38800
rect 1124 38548 1176 38554
rect 1124 38490 1176 38496
rect 1032 37256 1084 37262
rect 1032 37198 1084 37204
rect 1044 31090 1072 37198
rect 1136 36242 1164 38490
rect 1216 36712 1268 36718
rect 1216 36654 1268 36660
rect 1124 36236 1176 36242
rect 1124 36178 1176 36184
rect 1044 31062 1164 31090
rect 940 27600 992 27606
rect 940 27542 992 27548
rect 848 27056 900 27062
rect 848 26998 900 27004
rect 768 26206 1072 26234
rect 1044 21146 1072 26206
rect 1136 22098 1164 31062
rect 1228 24410 1256 36654
rect 1320 29714 1348 47602
rect 1412 32910 1440 49574
rect 1504 49230 1532 49642
rect 1492 49224 1544 49230
rect 1492 49166 1544 49172
rect 1492 49088 1544 49094
rect 1596 49076 1624 49778
rect 1544 49048 1624 49076
rect 1492 49030 1544 49036
rect 1492 48544 1544 48550
rect 1492 48486 1544 48492
rect 1504 48385 1532 48486
rect 1490 48376 1546 48385
rect 1490 48311 1546 48320
rect 1584 48340 1636 48346
rect 1584 48282 1636 48288
rect 1492 48000 1544 48006
rect 1492 47942 1544 47948
rect 1504 47841 1532 47942
rect 1490 47832 1546 47841
rect 1490 47767 1546 47776
rect 1492 47592 1544 47598
rect 1490 47560 1492 47569
rect 1544 47560 1546 47569
rect 1490 47495 1546 47504
rect 1492 47456 1544 47462
rect 1492 47398 1544 47404
rect 1504 47025 1532 47398
rect 1490 47016 1546 47025
rect 1490 46951 1546 46960
rect 1492 46912 1544 46918
rect 1492 46854 1544 46860
rect 1504 46617 1532 46854
rect 1490 46608 1546 46617
rect 1490 46543 1546 46552
rect 1492 46368 1544 46374
rect 1492 46310 1544 46316
rect 1504 46209 1532 46310
rect 1490 46200 1546 46209
rect 1490 46135 1546 46144
rect 1596 45937 1624 48282
rect 1582 45928 1638 45937
rect 1582 45863 1638 45872
rect 1492 45824 1544 45830
rect 1490 45792 1492 45801
rect 1544 45792 1546 45801
rect 1688 45778 1716 50118
rect 1490 45727 1546 45736
rect 1596 45750 1716 45778
rect 1492 45280 1544 45286
rect 1492 45222 1544 45228
rect 1504 45082 1532 45222
rect 1492 45076 1544 45082
rect 1492 45018 1544 45024
rect 1490 44840 1546 44849
rect 1490 44775 1546 44784
rect 1504 44538 1532 44775
rect 1492 44532 1544 44538
rect 1492 44474 1544 44480
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1504 41449 1532 41958
rect 1490 41440 1546 41449
rect 1490 41375 1546 41384
rect 1492 40384 1544 40390
rect 1492 40326 1544 40332
rect 1504 39681 1532 40326
rect 1490 39672 1546 39681
rect 1490 39607 1546 39616
rect 1492 39432 1544 39438
rect 1492 39374 1544 39380
rect 1504 38418 1532 39374
rect 1492 38412 1544 38418
rect 1492 38354 1544 38360
rect 1492 38208 1544 38214
rect 1492 38150 1544 38156
rect 1504 37777 1532 38150
rect 1490 37768 1546 37777
rect 1490 37703 1546 37712
rect 1492 37664 1544 37670
rect 1492 37606 1544 37612
rect 1504 37097 1532 37606
rect 1490 37088 1546 37097
rect 1490 37023 1546 37032
rect 1492 36576 1544 36582
rect 1492 36518 1544 36524
rect 1504 35873 1532 36518
rect 1490 35864 1546 35873
rect 1490 35799 1546 35808
rect 1490 35048 1546 35057
rect 1490 34983 1546 34992
rect 1504 34202 1532 34983
rect 1492 34196 1544 34202
rect 1492 34138 1544 34144
rect 1596 33522 1624 45750
rect 1676 45620 1728 45626
rect 1676 45562 1728 45568
rect 1688 43790 1716 45562
rect 1780 45014 1808 52006
rect 1872 45286 1900 52430
rect 1964 52154 1992 52550
rect 1952 52148 2004 52154
rect 1952 52090 2004 52096
rect 1952 50516 2004 50522
rect 1952 50458 2004 50464
rect 1964 50318 1992 50458
rect 1952 50312 2004 50318
rect 1952 50254 2004 50260
rect 1964 49842 1992 50254
rect 1952 49836 2004 49842
rect 1952 49778 2004 49784
rect 1952 49632 2004 49638
rect 1952 49574 2004 49580
rect 1964 48385 1992 49574
rect 1950 48376 2006 48385
rect 1950 48311 2006 48320
rect 1952 48136 2004 48142
rect 1952 48078 2004 48084
rect 1964 47190 1992 48078
rect 1952 47184 2004 47190
rect 1952 47126 2004 47132
rect 1952 46572 2004 46578
rect 1952 46514 2004 46520
rect 1964 45626 1992 46514
rect 1952 45620 2004 45626
rect 1952 45562 2004 45568
rect 1952 45484 2004 45490
rect 1952 45426 2004 45432
rect 1860 45280 1912 45286
rect 1860 45222 1912 45228
rect 1858 45112 1914 45121
rect 1858 45047 1914 45056
rect 1768 45008 1820 45014
rect 1768 44950 1820 44956
rect 1768 44396 1820 44402
rect 1768 44338 1820 44344
rect 1676 43784 1728 43790
rect 1676 43726 1728 43732
rect 1688 42786 1716 43726
rect 1780 42888 1808 44338
rect 1872 43790 1900 45047
rect 1860 43784 1912 43790
rect 1860 43726 1912 43732
rect 1780 42860 1900 42888
rect 1688 42758 1808 42786
rect 1676 42628 1728 42634
rect 1676 42570 1728 42576
rect 1688 42090 1716 42570
rect 1676 42084 1728 42090
rect 1676 42026 1728 42032
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1492 33312 1544 33318
rect 1492 33254 1544 33260
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1504 32473 1532 33254
rect 1688 32774 1716 42026
rect 1780 41614 1808 42758
rect 1872 41750 1900 42860
rect 1860 41744 1912 41750
rect 1860 41686 1912 41692
rect 1768 41608 1820 41614
rect 1768 41550 1820 41556
rect 1860 41608 1912 41614
rect 1860 41550 1912 41556
rect 1768 41472 1820 41478
rect 1768 41414 1820 41420
rect 1780 40526 1808 41414
rect 1768 40520 1820 40526
rect 1768 40462 1820 40468
rect 1872 40372 1900 41550
rect 1964 41290 1992 45426
rect 2056 41414 2084 55014
rect 2148 47530 2176 55916
rect 2332 55842 2360 57446
rect 2424 56982 2452 58006
rect 2412 56976 2464 56982
rect 2412 56918 2464 56924
rect 2412 56840 2464 56846
rect 2412 56782 2464 56788
rect 2240 55814 2360 55842
rect 2240 52698 2268 55814
rect 2320 55616 2372 55622
rect 2318 55584 2320 55593
rect 2372 55584 2374 55593
rect 2318 55519 2374 55528
rect 2320 55276 2372 55282
rect 2320 55218 2372 55224
rect 2332 54874 2360 55218
rect 2320 54868 2372 54874
rect 2320 54810 2372 54816
rect 2320 52896 2372 52902
rect 2320 52838 2372 52844
rect 2228 52692 2280 52698
rect 2228 52634 2280 52640
rect 2332 52601 2360 52838
rect 2318 52592 2374 52601
rect 2318 52527 2374 52536
rect 2320 52488 2372 52494
rect 2320 52430 2372 52436
rect 2228 51264 2280 51270
rect 2228 51206 2280 51212
rect 2240 50969 2268 51206
rect 2226 50960 2282 50969
rect 2226 50895 2282 50904
rect 2332 50674 2360 52430
rect 2240 50646 2360 50674
rect 2240 49280 2268 50646
rect 2424 50538 2452 56782
rect 2332 50510 2452 50538
rect 2516 50522 2544 60143
rect 2596 60104 2648 60110
rect 2596 60046 2648 60052
rect 2608 59634 2636 60046
rect 2686 59664 2742 59673
rect 2596 59628 2648 59634
rect 2686 59599 2688 59608
rect 2596 59570 2648 59576
rect 2740 59599 2742 59608
rect 2688 59570 2740 59576
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2596 57928 2648 57934
rect 2596 57870 2648 57876
rect 2608 57594 2636 57870
rect 2780 57792 2832 57798
rect 2778 57760 2780 57769
rect 2832 57760 2834 57769
rect 2778 57695 2834 57704
rect 2596 57588 2648 57594
rect 2596 57530 2648 57536
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2976 57050 3004 60706
rect 3054 59528 3110 59537
rect 3054 59463 3056 59472
rect 3108 59463 3110 59472
rect 3056 59434 3108 59440
rect 3056 57928 3108 57934
rect 3054 57896 3056 57905
rect 3108 57896 3110 57905
rect 3054 57831 3110 57840
rect 2964 57044 3016 57050
rect 2964 56986 3016 56992
rect 2596 56976 2648 56982
rect 2596 56918 2648 56924
rect 2608 56438 2636 56918
rect 2596 56432 2648 56438
rect 2596 56374 2648 56380
rect 2964 56432 3016 56438
rect 2964 56374 3016 56380
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2976 55962 3004 56374
rect 2964 55956 3016 55962
rect 2964 55898 3016 55904
rect 3056 55752 3108 55758
rect 3056 55694 3108 55700
rect 3068 55282 3096 55694
rect 3056 55276 3108 55282
rect 3056 55218 3108 55224
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 2780 54528 2832 54534
rect 2780 54470 2832 54476
rect 2792 54369 2820 54470
rect 2778 54360 2834 54369
rect 2778 54295 2834 54304
rect 2872 54188 2924 54194
rect 2872 54130 2924 54136
rect 2884 54074 2912 54130
rect 2884 54046 3004 54074
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2976 53514 3004 54046
rect 2596 53508 2648 53514
rect 2596 53450 2648 53456
rect 2964 53508 3016 53514
rect 2964 53450 3016 53456
rect 2608 52970 2636 53450
rect 3054 53000 3110 53009
rect 2596 52964 2648 52970
rect 3054 52935 3056 52944
rect 2596 52906 2648 52912
rect 3108 52935 3110 52944
rect 3056 52906 3108 52912
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2596 52556 2648 52562
rect 2596 52498 2648 52504
rect 2608 52018 2636 52498
rect 2596 52012 2648 52018
rect 2596 51954 2648 51960
rect 2964 52012 3016 52018
rect 2964 51954 3016 51960
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2780 51400 2832 51406
rect 2780 51342 2832 51348
rect 2792 50794 2820 51342
rect 2780 50788 2832 50794
rect 2780 50730 2832 50736
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2504 50516 2556 50522
rect 2332 49638 2360 50510
rect 2504 50458 2556 50464
rect 2412 50448 2464 50454
rect 2412 50390 2464 50396
rect 2424 49722 2452 50390
rect 2976 50318 3004 51954
rect 3054 51368 3110 51377
rect 3054 51303 3110 51312
rect 3068 51270 3096 51303
rect 3056 51264 3108 51270
rect 3056 51206 3108 51212
rect 2964 50312 3016 50318
rect 3016 50272 3096 50300
rect 2964 50254 3016 50260
rect 2424 49694 2544 49722
rect 2320 49632 2372 49638
rect 2412 49632 2464 49638
rect 2320 49574 2372 49580
rect 2410 49600 2412 49609
rect 2464 49600 2466 49609
rect 2410 49535 2466 49544
rect 2240 49252 2452 49280
rect 2226 49192 2282 49201
rect 2226 49127 2282 49136
rect 2240 48890 2268 49127
rect 2320 49088 2372 49094
rect 2320 49030 2372 49036
rect 2228 48884 2280 48890
rect 2228 48826 2280 48832
rect 2228 48612 2280 48618
rect 2228 48554 2280 48560
rect 2136 47524 2188 47530
rect 2136 47466 2188 47472
rect 2240 47274 2268 48554
rect 2148 47246 2268 47274
rect 2148 44266 2176 47246
rect 2228 47184 2280 47190
rect 2228 47126 2280 47132
rect 2240 45393 2268 47126
rect 2226 45384 2282 45393
rect 2226 45319 2282 45328
rect 2240 44946 2268 45319
rect 2228 44940 2280 44946
rect 2228 44882 2280 44888
rect 2332 44282 2360 49030
rect 2424 48618 2452 49252
rect 2412 48612 2464 48618
rect 2412 48554 2464 48560
rect 2412 48340 2464 48346
rect 2412 48282 2464 48288
rect 2424 44402 2452 48282
rect 2516 47734 2544 49694
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2780 49088 2832 49094
rect 2780 49030 2832 49036
rect 2792 48793 2820 49030
rect 2778 48784 2834 48793
rect 2778 48719 2834 48728
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2582 48368 2890 48388
rect 2962 48328 3018 48337
rect 2872 48272 2924 48278
rect 3068 48278 3096 50272
rect 2962 48263 3018 48272
rect 3056 48272 3108 48278
rect 2872 48214 2924 48220
rect 2780 48136 2832 48142
rect 2780 48078 2832 48084
rect 2792 47841 2820 48078
rect 2778 47832 2834 47841
rect 2778 47767 2834 47776
rect 2504 47728 2556 47734
rect 2504 47670 2556 47676
rect 2884 47666 2912 48214
rect 2976 47802 3004 48263
rect 3056 48214 3108 48220
rect 3056 48136 3108 48142
rect 3056 48078 3108 48084
rect 2964 47796 3016 47802
rect 2964 47738 3016 47744
rect 2688 47660 2740 47666
rect 2688 47602 2740 47608
rect 2872 47660 2924 47666
rect 2872 47602 2924 47608
rect 2964 47660 3016 47666
rect 2964 47602 3016 47608
rect 2504 47592 2556 47598
rect 2700 47569 2728 47602
rect 2504 47534 2556 47540
rect 2686 47560 2742 47569
rect 2516 47054 2544 47534
rect 2686 47495 2742 47504
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2504 47048 2556 47054
rect 2504 46990 2556 46996
rect 2872 47048 2924 47054
rect 2872 46990 2924 46996
rect 2516 45014 2544 46990
rect 2596 46912 2648 46918
rect 2596 46854 2648 46860
rect 2780 46912 2832 46918
rect 2780 46854 2832 46860
rect 2608 46646 2636 46854
rect 2596 46640 2648 46646
rect 2596 46582 2648 46588
rect 2792 46578 2820 46854
rect 2884 46714 2912 46990
rect 2872 46708 2924 46714
rect 2872 46650 2924 46656
rect 2780 46572 2832 46578
rect 2780 46514 2832 46520
rect 2792 46481 2820 46514
rect 2778 46472 2834 46481
rect 2778 46407 2834 46416
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2504 45008 2556 45014
rect 2780 45008 2832 45014
rect 2504 44950 2556 44956
rect 2778 44976 2780 44985
rect 2832 44976 2834 44985
rect 2412 44396 2464 44402
rect 2412 44338 2464 44344
rect 2136 44260 2188 44266
rect 2136 44202 2188 44208
rect 2240 44254 2360 44282
rect 2412 44260 2464 44266
rect 2136 43852 2188 43858
rect 2136 43794 2188 43800
rect 2148 43382 2176 43794
rect 2136 43376 2188 43382
rect 2136 43318 2188 43324
rect 2148 42702 2176 43318
rect 2136 42696 2188 42702
rect 2136 42638 2188 42644
rect 2148 41614 2176 42638
rect 2240 42106 2268 44254
rect 2412 44202 2464 44208
rect 2320 44192 2372 44198
rect 2320 44134 2372 44140
rect 2332 43625 2360 44134
rect 2318 43616 2374 43625
rect 2318 43551 2374 43560
rect 2424 42226 2452 44202
rect 2516 43858 2544 44950
rect 2778 44911 2834 44920
rect 2976 44826 3004 47602
rect 3068 47258 3096 48078
rect 3056 47252 3108 47258
rect 3056 47194 3108 47200
rect 2976 44798 3096 44826
rect 2780 44736 2832 44742
rect 2780 44678 2832 44684
rect 2792 44441 2820 44678
rect 2778 44432 2834 44441
rect 2778 44367 2834 44376
rect 2964 44192 3016 44198
rect 2964 44134 3016 44140
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2976 43897 3004 44134
rect 2962 43888 3018 43897
rect 2504 43852 2556 43858
rect 2962 43823 3018 43832
rect 2504 43794 2556 43800
rect 2964 43716 3016 43722
rect 2964 43658 3016 43664
rect 2780 43648 2832 43654
rect 2780 43590 2832 43596
rect 2792 43217 2820 43590
rect 2976 43382 3004 43658
rect 3068 43382 3096 44798
rect 3160 44402 3188 60998
rect 3252 60734 3280 66574
rect 3332 65408 3384 65414
rect 3332 65350 3384 65356
rect 3344 65113 3372 65350
rect 3330 65104 3386 65113
rect 3330 65039 3386 65048
rect 3424 65068 3476 65074
rect 3424 65010 3476 65016
rect 3436 64954 3464 65010
rect 3344 64926 3464 64954
rect 3344 62898 3372 64926
rect 3424 64864 3476 64870
rect 3424 64806 3476 64812
rect 3332 62892 3384 62898
rect 3332 62834 3384 62840
rect 3344 61198 3372 62834
rect 3332 61192 3384 61198
rect 3332 61134 3384 61140
rect 3252 60706 3372 60734
rect 3240 59424 3292 59430
rect 3240 59366 3292 59372
rect 3252 57798 3280 59366
rect 3240 57792 3292 57798
rect 3240 57734 3292 57740
rect 3344 57594 3372 60706
rect 3332 57588 3384 57594
rect 3332 57530 3384 57536
rect 3240 57452 3292 57458
rect 3240 57394 3292 57400
rect 3252 56370 3280 57394
rect 3332 57384 3384 57390
rect 3332 57326 3384 57332
rect 3344 56846 3372 57326
rect 3332 56840 3384 56846
rect 3332 56782 3384 56788
rect 3240 56364 3292 56370
rect 3240 56306 3292 56312
rect 3240 56228 3292 56234
rect 3240 56170 3292 56176
rect 3148 44396 3200 44402
rect 3148 44338 3200 44344
rect 3252 44282 3280 56170
rect 3344 55350 3372 56782
rect 3332 55344 3384 55350
rect 3332 55286 3384 55292
rect 3344 53582 3372 55286
rect 3332 53576 3384 53582
rect 3332 53518 3384 53524
rect 3344 52562 3372 53518
rect 3332 52556 3384 52562
rect 3332 52498 3384 52504
rect 3332 51876 3384 51882
rect 3332 51818 3384 51824
rect 3160 44254 3280 44282
rect 2964 43376 3016 43382
rect 2964 43318 3016 43324
rect 3056 43376 3108 43382
rect 3056 43318 3108 43324
rect 2778 43208 2834 43217
rect 2778 43143 2834 43152
rect 2964 43104 3016 43110
rect 2964 43046 3016 43052
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2872 42832 2924 42838
rect 2872 42774 2924 42780
rect 2504 42628 2556 42634
rect 2504 42570 2556 42576
rect 2412 42220 2464 42226
rect 2412 42162 2464 42168
rect 2240 42078 2452 42106
rect 2228 42016 2280 42022
rect 2228 41958 2280 41964
rect 2240 41857 2268 41958
rect 2226 41848 2282 41857
rect 2226 41783 2282 41792
rect 2228 41676 2280 41682
rect 2280 41636 2360 41664
rect 2228 41618 2280 41624
rect 2136 41608 2188 41614
rect 2136 41550 2188 41556
rect 2056 41386 2268 41414
rect 1964 41262 2176 41290
rect 2044 41064 2096 41070
rect 2044 41006 2096 41012
rect 1950 40896 2006 40905
rect 1950 40831 2006 40840
rect 1780 40344 1900 40372
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 1676 32768 1728 32774
rect 1676 32710 1728 32716
rect 1490 32464 1546 32473
rect 1490 32399 1546 32408
rect 1492 32224 1544 32230
rect 1492 32166 1544 32172
rect 1504 31113 1532 32166
rect 1596 31929 1624 32710
rect 1780 32586 1808 40344
rect 1860 40180 1912 40186
rect 1860 40122 1912 40128
rect 1872 40050 1900 40122
rect 1860 40044 1912 40050
rect 1860 39986 1912 39992
rect 1872 39438 1900 39986
rect 1860 39432 1912 39438
rect 1860 39374 1912 39380
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 1688 32558 1808 32586
rect 1582 31920 1638 31929
rect 1582 31855 1638 31864
rect 1490 31104 1546 31113
rect 1688 31090 1716 32558
rect 1768 32360 1820 32366
rect 1768 32302 1820 32308
rect 1490 31039 1546 31048
rect 1596 31062 1716 31090
rect 1490 30696 1546 30705
rect 1490 30631 1546 30640
rect 1504 30122 1532 30631
rect 1492 30116 1544 30122
rect 1492 30058 1544 30064
rect 1596 30002 1624 31062
rect 1676 30864 1728 30870
rect 1676 30806 1728 30812
rect 1688 30258 1716 30806
rect 1676 30252 1728 30258
rect 1676 30194 1728 30200
rect 1780 30138 1808 32302
rect 1872 31929 1900 38898
rect 1964 32910 1992 40831
rect 2056 33522 2084 41006
rect 2148 40168 2176 41262
rect 2240 41070 2268 41386
rect 2228 41064 2280 41070
rect 2228 41006 2280 41012
rect 2228 40928 2280 40934
rect 2228 40870 2280 40876
rect 2240 40633 2268 40870
rect 2226 40624 2282 40633
rect 2226 40559 2282 40568
rect 2148 40140 2268 40168
rect 2134 40080 2190 40089
rect 2134 40015 2190 40024
rect 2148 38418 2176 40015
rect 2240 39930 2268 40140
rect 2332 40050 2360 41636
rect 2424 41596 2452 42078
rect 2516 41698 2544 42570
rect 2884 42276 2912 42774
rect 2976 42673 3004 43046
rect 2962 42664 3018 42673
rect 2962 42599 3018 42608
rect 3056 42560 3108 42566
rect 3056 42502 3108 42508
rect 2964 42288 3016 42294
rect 2884 42248 2964 42276
rect 3068 42265 3096 42502
rect 2964 42230 3016 42236
rect 3054 42256 3110 42265
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2516 41670 2636 41698
rect 2424 41568 2544 41596
rect 2412 41472 2464 41478
rect 2412 41414 2464 41420
rect 2320 40044 2372 40050
rect 2320 39986 2372 39992
rect 2240 39902 2360 39930
rect 2228 39840 2280 39846
rect 2228 39782 2280 39788
rect 2136 38412 2188 38418
rect 2136 38354 2188 38360
rect 2136 38276 2188 38282
rect 2136 38218 2188 38224
rect 2148 37874 2176 38218
rect 2136 37868 2188 37874
rect 2136 37810 2188 37816
rect 2148 37398 2176 37810
rect 2136 37392 2188 37398
rect 2136 37334 2188 37340
rect 2240 37097 2268 39782
rect 2226 37088 2282 37097
rect 2226 37023 2282 37032
rect 2332 36854 2360 39902
rect 2320 36848 2372 36854
rect 2226 36816 2282 36825
rect 2320 36790 2372 36796
rect 2226 36751 2282 36760
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 2148 34610 2176 35022
rect 2136 34604 2188 34610
rect 2136 34546 2188 34552
rect 2136 34468 2188 34474
rect 2136 34410 2188 34416
rect 2148 33998 2176 34410
rect 2136 33992 2188 33998
rect 2136 33934 2188 33940
rect 2044 33516 2096 33522
rect 2044 33458 2096 33464
rect 2136 33380 2188 33386
rect 2136 33322 2188 33328
rect 1952 32904 2004 32910
rect 1952 32846 2004 32852
rect 1952 32768 2004 32774
rect 1952 32710 2004 32716
rect 1858 31920 1914 31929
rect 1858 31855 1914 31864
rect 1858 31784 1914 31793
rect 1858 31719 1914 31728
rect 1504 29974 1624 30002
rect 1688 30110 1808 30138
rect 1308 29708 1360 29714
rect 1308 29650 1360 29656
rect 1308 29232 1360 29238
rect 1308 29174 1360 29180
rect 1216 24404 1268 24410
rect 1216 24346 1268 24352
rect 1216 23724 1268 23730
rect 1216 23666 1268 23672
rect 1228 22137 1256 23666
rect 1214 22128 1270 22137
rect 1124 22092 1176 22098
rect 1214 22063 1270 22072
rect 1124 22034 1176 22040
rect 1032 21140 1084 21146
rect 1032 21082 1084 21088
rect 1320 17218 1348 29174
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28121 1440 29106
rect 1398 28112 1454 28121
rect 1398 28047 1454 28056
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 26353 1440 27406
rect 1504 26586 1532 29974
rect 1584 29640 1636 29646
rect 1584 29582 1636 29588
rect 1596 29306 1624 29582
rect 1584 29300 1636 29306
rect 1584 29242 1636 29248
rect 1584 29164 1636 29170
rect 1584 29106 1636 29112
rect 1492 26580 1544 26586
rect 1492 26522 1544 26528
rect 1398 26344 1454 26353
rect 1398 26279 1454 26288
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1492 25900 1544 25906
rect 1492 25842 1544 25848
rect 1412 24313 1440 25842
rect 1504 25129 1532 25842
rect 1490 25120 1546 25129
rect 1490 25055 1546 25064
rect 1492 24812 1544 24818
rect 1492 24754 1544 24760
rect 1398 24304 1454 24313
rect 1398 24239 1454 24248
rect 1400 23520 1452 23526
rect 1400 23462 1452 23468
rect 1412 22642 1440 23462
rect 1504 22953 1532 24754
rect 1490 22944 1546 22953
rect 1490 22879 1546 22888
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1492 21616 1544 21622
rect 1492 21558 1544 21564
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21185 1440 21490
rect 1398 21176 1454 21185
rect 1398 21111 1454 21120
rect 1504 17354 1532 21558
rect 1596 17814 1624 29106
rect 1688 28218 1716 30110
rect 1768 29572 1820 29578
rect 1768 29514 1820 29520
rect 1780 29102 1808 29514
rect 1768 29096 1820 29102
rect 1768 29038 1820 29044
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1780 28218 1808 28494
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 1768 28212 1820 28218
rect 1768 28154 1820 28160
rect 1766 28112 1822 28121
rect 1766 28047 1822 28056
rect 1676 27940 1728 27946
rect 1676 27882 1728 27888
rect 1688 26234 1716 27882
rect 1780 26382 1808 28047
rect 1872 26858 1900 31719
rect 1860 26852 1912 26858
rect 1860 26794 1912 26800
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1688 26206 1808 26234
rect 1676 24268 1728 24274
rect 1676 24210 1728 24216
rect 1688 23118 1716 24210
rect 1676 23112 1728 23118
rect 1676 23054 1728 23060
rect 1688 18426 1716 23054
rect 1780 18970 1808 26206
rect 1964 24750 1992 32710
rect 2044 32428 2096 32434
rect 2044 32370 2096 32376
rect 2056 27946 2084 32370
rect 2148 31142 2176 33322
rect 2240 32586 2268 36751
rect 2320 36576 2372 36582
rect 2320 36518 2372 36524
rect 2332 36281 2360 36518
rect 2318 36272 2374 36281
rect 2318 36207 2374 36216
rect 2320 35692 2372 35698
rect 2320 35634 2372 35640
rect 2332 33946 2360 35634
rect 2424 34610 2452 41414
rect 2412 34604 2464 34610
rect 2412 34546 2464 34552
rect 2412 34400 2464 34406
rect 2412 34342 2464 34348
rect 2424 34105 2452 34342
rect 2516 34184 2544 41568
rect 2608 41177 2636 41670
rect 2688 41676 2740 41682
rect 2688 41618 2740 41624
rect 2594 41168 2650 41177
rect 2700 41138 2728 41618
rect 2976 41614 3004 42230
rect 3054 42191 3110 42200
rect 2964 41608 3016 41614
rect 2964 41550 3016 41556
rect 2594 41103 2650 41112
rect 2688 41132 2740 41138
rect 2688 41074 2740 41080
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2872 40520 2924 40526
rect 2872 40462 2924 40468
rect 2596 40452 2648 40458
rect 2596 40394 2648 40400
rect 2608 40186 2636 40394
rect 2596 40180 2648 40186
rect 2596 40122 2648 40128
rect 2884 40050 2912 40462
rect 2872 40044 2924 40050
rect 2976 40032 3004 41550
rect 3054 41032 3110 41041
rect 3054 40967 3056 40976
rect 3108 40967 3110 40976
rect 3056 40938 3108 40944
rect 3056 40044 3108 40050
rect 2976 40004 3056 40032
rect 2872 39986 2924 39992
rect 3056 39986 3108 39992
rect 2884 39930 2912 39986
rect 2884 39902 3004 39930
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2872 39364 2924 39370
rect 2872 39306 2924 39312
rect 2780 39296 2832 39302
rect 2778 39264 2780 39273
rect 2832 39264 2834 39273
rect 2778 39199 2834 39208
rect 2884 38826 2912 39306
rect 2976 38894 3004 39902
rect 2964 38888 3016 38894
rect 2964 38830 3016 38836
rect 2872 38820 2924 38826
rect 2872 38762 2924 38768
rect 2964 38752 3016 38758
rect 2964 38694 3016 38700
rect 2582 38652 2890 38672
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2976 38049 3004 38694
rect 3068 38350 3096 39986
rect 3056 38344 3108 38350
rect 3056 38286 3108 38292
rect 2962 38040 3018 38049
rect 2962 37975 3018 37984
rect 2964 37868 3016 37874
rect 2964 37810 3016 37816
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2976 37398 3004 37810
rect 2964 37392 3016 37398
rect 2964 37334 3016 37340
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2976 36038 3004 37334
rect 3068 37262 3096 38286
rect 3056 37256 3108 37262
rect 3056 37198 3108 37204
rect 3054 36680 3110 36689
rect 3054 36615 3056 36624
rect 3108 36615 3110 36624
rect 3056 36586 3108 36592
rect 2964 36032 3016 36038
rect 2964 35974 3016 35980
rect 2976 35630 3004 35974
rect 2964 35624 3016 35630
rect 2964 35566 3016 35572
rect 3054 35592 3110 35601
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2976 35086 3004 35566
rect 3054 35527 3056 35536
rect 3108 35527 3110 35536
rect 3056 35498 3108 35504
rect 2964 35080 3016 35086
rect 2964 35022 3016 35028
rect 2964 34944 3016 34950
rect 2964 34886 3016 34892
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2516 34156 2636 34184
rect 2410 34096 2466 34105
rect 2410 34031 2466 34040
rect 2332 33918 2452 33946
rect 2320 33856 2372 33862
rect 2320 33798 2372 33804
rect 2332 33697 2360 33798
rect 2318 33688 2374 33697
rect 2318 33623 2374 33632
rect 2320 33312 2372 33318
rect 2318 33280 2320 33289
rect 2372 33280 2374 33289
rect 2318 33215 2374 33224
rect 2318 32872 2374 32881
rect 2318 32807 2374 32816
rect 2332 32774 2360 32807
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2240 32558 2360 32586
rect 2136 31136 2188 31142
rect 2136 31078 2188 31084
rect 2228 30252 2280 30258
rect 2228 30194 2280 30200
rect 2136 30184 2188 30190
rect 2136 30126 2188 30132
rect 2148 29782 2176 30126
rect 2136 29776 2188 29782
rect 2136 29718 2188 29724
rect 2148 29170 2176 29718
rect 2136 29164 2188 29170
rect 2136 29106 2188 29112
rect 2136 29028 2188 29034
rect 2136 28970 2188 28976
rect 2044 27940 2096 27946
rect 2044 27882 2096 27888
rect 2042 27568 2098 27577
rect 2042 27503 2098 27512
rect 1952 24744 2004 24750
rect 1952 24686 2004 24692
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1872 19378 1900 19654
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1860 18148 1912 18154
rect 1860 18090 1912 18096
rect 1584 17808 1636 17814
rect 1584 17750 1636 17756
rect 1504 17326 1716 17354
rect 1228 17190 1348 17218
rect 1400 17196 1452 17202
rect 1228 7478 1256 17190
rect 1400 17138 1452 17144
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1412 15609 1440 17138
rect 1504 16561 1532 17138
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1490 16552 1546 16561
rect 1490 16487 1546 16496
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1398 15600 1454 15609
rect 1398 15535 1454 15544
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1412 13410 1440 15098
rect 1504 14618 1532 16050
rect 1596 15502 1624 16934
rect 1688 16182 1716 17326
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1676 16176 1728 16182
rect 1676 16118 1728 16124
rect 1688 15994 1716 16118
rect 1780 16114 1808 16934
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1688 15966 1808 15994
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15706 1716 15846
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1584 15496 1636 15502
rect 1780 15450 1808 15966
rect 1584 15438 1636 15444
rect 1688 15422 1808 15450
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15094 1624 15302
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 14074 1532 14418
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1412 13382 1532 13410
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1320 11801 1348 12718
rect 1412 12345 1440 13262
rect 1504 12986 1532 13382
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1596 12434 1624 15030
rect 1688 14550 1716 15422
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1676 14544 1728 14550
rect 1676 14486 1728 14492
rect 1780 14482 1808 15302
rect 1872 15026 1900 18090
rect 1964 17882 1992 23666
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 2056 17218 2084 27503
rect 2148 27418 2176 28970
rect 2240 27554 2268 30194
rect 2332 28762 2360 32558
rect 2424 32434 2452 33918
rect 2608 33674 2636 34156
rect 2516 33646 2636 33674
rect 2412 32428 2464 32434
rect 2412 32370 2464 32376
rect 2516 31822 2544 33646
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2976 32910 3004 34886
rect 3056 34740 3108 34746
rect 3056 34682 3108 34688
rect 3068 33862 3096 34682
rect 3160 34610 3188 44254
rect 3240 44192 3292 44198
rect 3240 44134 3292 44140
rect 3252 38962 3280 44134
rect 3344 41274 3372 51818
rect 3436 45558 3464 64806
rect 3528 59974 3556 69158
rect 3620 64870 3648 69974
rect 3792 66768 3844 66774
rect 3792 66710 3844 66716
rect 3608 64864 3660 64870
rect 3608 64806 3660 64812
rect 3700 63980 3752 63986
rect 3700 63922 3752 63928
rect 3608 61328 3660 61334
rect 3608 61270 3660 61276
rect 3516 59968 3568 59974
rect 3516 59910 3568 59916
rect 3516 58064 3568 58070
rect 3516 58006 3568 58012
rect 3528 56953 3556 58006
rect 3514 56944 3570 56953
rect 3514 56879 3570 56888
rect 3516 56772 3568 56778
rect 3516 56714 3568 56720
rect 3528 56370 3556 56714
rect 3620 56438 3648 61270
rect 3608 56432 3660 56438
rect 3608 56374 3660 56380
rect 3516 56364 3568 56370
rect 3516 56306 3568 56312
rect 3528 54194 3556 56306
rect 3608 54800 3660 54806
rect 3608 54742 3660 54748
rect 3516 54188 3568 54194
rect 3516 54130 3568 54136
rect 3528 52018 3556 54130
rect 3516 52012 3568 52018
rect 3516 51954 3568 51960
rect 3528 50998 3556 51954
rect 3516 50992 3568 50998
rect 3516 50934 3568 50940
rect 3528 50454 3556 50934
rect 3516 50448 3568 50454
rect 3516 50390 3568 50396
rect 3528 49230 3556 50390
rect 3516 49224 3568 49230
rect 3516 49166 3568 49172
rect 3516 49088 3568 49094
rect 3516 49030 3568 49036
rect 3528 47841 3556 49030
rect 3514 47832 3570 47841
rect 3514 47767 3516 47776
rect 3568 47767 3570 47776
rect 3516 47738 3568 47744
rect 3516 47660 3568 47666
rect 3516 47602 3568 47608
rect 3528 47190 3556 47602
rect 3516 47184 3568 47190
rect 3516 47126 3568 47132
rect 3620 47002 3648 54742
rect 3712 50522 3740 63922
rect 3804 61266 3832 66710
rect 3884 64932 3936 64938
rect 3884 64874 3936 64880
rect 3896 64569 3924 64874
rect 3882 64560 3938 64569
rect 3882 64495 3938 64504
rect 3792 61260 3844 61266
rect 3792 61202 3844 61208
rect 3884 61192 3936 61198
rect 3884 61134 3936 61140
rect 3792 59016 3844 59022
rect 3792 58958 3844 58964
rect 3804 51074 3832 58958
rect 3896 57934 3924 61134
rect 3884 57928 3936 57934
rect 3884 57870 3936 57876
rect 3884 57792 3936 57798
rect 3884 57734 3936 57740
rect 3896 56234 3924 57734
rect 3884 56228 3936 56234
rect 3884 56170 3936 56176
rect 3804 51046 3924 51074
rect 3792 50788 3844 50794
rect 3792 50730 3844 50736
rect 3700 50516 3752 50522
rect 3700 50458 3752 50464
rect 3698 50416 3754 50425
rect 3698 50351 3754 50360
rect 3712 47161 3740 50351
rect 3698 47152 3754 47161
rect 3698 47087 3754 47096
rect 3620 46974 3740 47002
rect 3516 46572 3568 46578
rect 3516 46514 3568 46520
rect 3424 45552 3476 45558
rect 3424 45494 3476 45500
rect 3422 45384 3478 45393
rect 3422 45319 3478 45328
rect 3436 41585 3464 45319
rect 3422 41576 3478 41585
rect 3422 41511 3478 41520
rect 3424 41472 3476 41478
rect 3424 41414 3476 41420
rect 3332 41268 3384 41274
rect 3332 41210 3384 41216
rect 3330 41168 3386 41177
rect 3330 41103 3386 41112
rect 3240 38956 3292 38962
rect 3240 38898 3292 38904
rect 3240 38820 3292 38826
rect 3240 38762 3292 38768
rect 3252 37369 3280 38762
rect 3238 37360 3294 37369
rect 3238 37295 3294 37304
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 3252 36378 3280 37198
rect 3240 36372 3292 36378
rect 3240 36314 3292 36320
rect 3240 34740 3292 34746
rect 3240 34682 3292 34688
rect 3148 34604 3200 34610
rect 3148 34546 3200 34552
rect 3252 34513 3280 34682
rect 3238 34504 3294 34513
rect 3238 34439 3294 34448
rect 3344 34354 3372 41103
rect 3436 39438 3464 41414
rect 3424 39432 3476 39438
rect 3424 39374 3476 39380
rect 3528 39098 3556 46514
rect 3712 46322 3740 46974
rect 3804 46578 3832 50730
rect 3792 46572 3844 46578
rect 3792 46514 3844 46520
rect 3712 46294 3832 46322
rect 3608 46096 3660 46102
rect 3608 46038 3660 46044
rect 3620 43976 3648 46038
rect 3804 44198 3832 46294
rect 3792 44192 3844 44198
rect 3792 44134 3844 44140
rect 3620 43948 3740 43976
rect 3608 43784 3660 43790
rect 3608 43726 3660 43732
rect 3620 43314 3648 43726
rect 3608 43308 3660 43314
rect 3608 43250 3660 43256
rect 3608 43172 3660 43178
rect 3608 43114 3660 43120
rect 3620 41546 3648 43114
rect 3712 42702 3740 43948
rect 3896 43450 3924 51046
rect 3988 49858 4016 75686
rect 4213 75100 4521 75120
rect 4213 75098 4219 75100
rect 4275 75098 4299 75100
rect 4355 75098 4379 75100
rect 4435 75098 4459 75100
rect 4515 75098 4521 75100
rect 4275 75046 4277 75098
rect 4457 75046 4459 75098
rect 4213 75044 4219 75046
rect 4275 75044 4299 75046
rect 4355 75044 4379 75046
rect 4435 75044 4459 75046
rect 4515 75044 4521 75046
rect 4213 75024 4521 75044
rect 4213 74012 4521 74032
rect 4213 74010 4219 74012
rect 4275 74010 4299 74012
rect 4355 74010 4379 74012
rect 4435 74010 4459 74012
rect 4515 74010 4521 74012
rect 4275 73958 4277 74010
rect 4457 73958 4459 74010
rect 4213 73956 4219 73958
rect 4275 73956 4299 73958
rect 4355 73956 4379 73958
rect 4435 73956 4459 73958
rect 4515 73956 4521 73958
rect 4213 73936 4521 73956
rect 4068 73092 4120 73098
rect 4068 73034 4120 73040
rect 4080 72622 4108 73034
rect 4213 72924 4521 72944
rect 4213 72922 4219 72924
rect 4275 72922 4299 72924
rect 4355 72922 4379 72924
rect 4435 72922 4459 72924
rect 4515 72922 4521 72924
rect 4275 72870 4277 72922
rect 4457 72870 4459 72922
rect 4213 72868 4219 72870
rect 4275 72868 4299 72870
rect 4355 72868 4379 72870
rect 4435 72868 4459 72870
rect 4515 72868 4521 72870
rect 4213 72848 4521 72868
rect 4068 72616 4120 72622
rect 4068 72558 4120 72564
rect 4213 71836 4521 71856
rect 4213 71834 4219 71836
rect 4275 71834 4299 71836
rect 4355 71834 4379 71836
rect 4435 71834 4459 71836
rect 4515 71834 4521 71836
rect 4275 71782 4277 71834
rect 4457 71782 4459 71834
rect 4213 71780 4219 71782
rect 4275 71780 4299 71782
rect 4355 71780 4379 71782
rect 4435 71780 4459 71782
rect 4515 71780 4521 71782
rect 4213 71760 4521 71780
rect 5080 71120 5132 71126
rect 5080 71062 5132 71068
rect 4213 70748 4521 70768
rect 4213 70746 4219 70748
rect 4275 70746 4299 70748
rect 4355 70746 4379 70748
rect 4435 70746 4459 70748
rect 4515 70746 4521 70748
rect 4275 70694 4277 70746
rect 4457 70694 4459 70746
rect 4213 70692 4219 70694
rect 4275 70692 4299 70694
rect 4355 70692 4379 70694
rect 4435 70692 4459 70694
rect 4515 70692 4521 70694
rect 4213 70672 4521 70692
rect 4213 69660 4521 69680
rect 4213 69658 4219 69660
rect 4275 69658 4299 69660
rect 4355 69658 4379 69660
rect 4435 69658 4459 69660
rect 4515 69658 4521 69660
rect 4275 69606 4277 69658
rect 4457 69606 4459 69658
rect 4213 69604 4219 69606
rect 4275 69604 4299 69606
rect 4355 69604 4379 69606
rect 4435 69604 4459 69606
rect 4515 69604 4521 69606
rect 4213 69584 4521 69604
rect 4213 68572 4521 68592
rect 4213 68570 4219 68572
rect 4275 68570 4299 68572
rect 4355 68570 4379 68572
rect 4435 68570 4459 68572
rect 4515 68570 4521 68572
rect 4275 68518 4277 68570
rect 4457 68518 4459 68570
rect 4213 68516 4219 68518
rect 4275 68516 4299 68518
rect 4355 68516 4379 68518
rect 4435 68516 4459 68518
rect 4515 68516 4521 68518
rect 4213 68496 4521 68516
rect 4213 67484 4521 67504
rect 4213 67482 4219 67484
rect 4275 67482 4299 67484
rect 4355 67482 4379 67484
rect 4435 67482 4459 67484
rect 4515 67482 4521 67484
rect 4275 67430 4277 67482
rect 4457 67430 4459 67482
rect 4213 67428 4219 67430
rect 4275 67428 4299 67430
rect 4355 67428 4379 67430
rect 4435 67428 4459 67430
rect 4515 67428 4521 67430
rect 4213 67408 4521 67428
rect 4213 66396 4521 66416
rect 4213 66394 4219 66396
rect 4275 66394 4299 66396
rect 4355 66394 4379 66396
rect 4435 66394 4459 66396
rect 4515 66394 4521 66396
rect 4275 66342 4277 66394
rect 4457 66342 4459 66394
rect 4213 66340 4219 66342
rect 4275 66340 4299 66342
rect 4355 66340 4379 66342
rect 4435 66340 4459 66342
rect 4515 66340 4521 66342
rect 4213 66320 4521 66340
rect 4213 65308 4521 65328
rect 4213 65306 4219 65308
rect 4275 65306 4299 65308
rect 4355 65306 4379 65308
rect 4435 65306 4459 65308
rect 4515 65306 4521 65308
rect 4275 65254 4277 65306
rect 4457 65254 4459 65306
rect 4213 65252 4219 65254
rect 4275 65252 4299 65254
rect 4355 65252 4379 65254
rect 4435 65252 4459 65254
rect 4515 65252 4521 65254
rect 4213 65232 4521 65252
rect 4213 64220 4521 64240
rect 4213 64218 4219 64220
rect 4275 64218 4299 64220
rect 4355 64218 4379 64220
rect 4435 64218 4459 64220
rect 4515 64218 4521 64220
rect 4275 64166 4277 64218
rect 4457 64166 4459 64218
rect 4213 64164 4219 64166
rect 4275 64164 4299 64166
rect 4355 64164 4379 64166
rect 4435 64164 4459 64166
rect 4515 64164 4521 64166
rect 4213 64144 4521 64164
rect 4620 63912 4672 63918
rect 4620 63854 4672 63860
rect 4213 63132 4521 63152
rect 4213 63130 4219 63132
rect 4275 63130 4299 63132
rect 4355 63130 4379 63132
rect 4435 63130 4459 63132
rect 4515 63130 4521 63132
rect 4275 63078 4277 63130
rect 4457 63078 4459 63130
rect 4213 63076 4219 63078
rect 4275 63076 4299 63078
rect 4355 63076 4379 63078
rect 4435 63076 4459 63078
rect 4515 63076 4521 63078
rect 4213 63056 4521 63076
rect 4213 62044 4521 62064
rect 4213 62042 4219 62044
rect 4275 62042 4299 62044
rect 4355 62042 4379 62044
rect 4435 62042 4459 62044
rect 4515 62042 4521 62044
rect 4275 61990 4277 62042
rect 4457 61990 4459 62042
rect 4213 61988 4219 61990
rect 4275 61988 4299 61990
rect 4355 61988 4379 61990
rect 4435 61988 4459 61990
rect 4515 61988 4521 61990
rect 4213 61968 4521 61988
rect 4068 61396 4120 61402
rect 4068 61338 4120 61344
rect 4080 58070 4108 61338
rect 4213 60956 4521 60976
rect 4213 60954 4219 60956
rect 4275 60954 4299 60956
rect 4355 60954 4379 60956
rect 4435 60954 4459 60956
rect 4515 60954 4521 60956
rect 4275 60902 4277 60954
rect 4457 60902 4459 60954
rect 4213 60900 4219 60902
rect 4275 60900 4299 60902
rect 4355 60900 4379 60902
rect 4435 60900 4459 60902
rect 4515 60900 4521 60902
rect 4213 60880 4521 60900
rect 4213 59868 4521 59888
rect 4213 59866 4219 59868
rect 4275 59866 4299 59868
rect 4355 59866 4379 59868
rect 4435 59866 4459 59868
rect 4515 59866 4521 59868
rect 4275 59814 4277 59866
rect 4457 59814 4459 59866
rect 4213 59812 4219 59814
rect 4275 59812 4299 59814
rect 4355 59812 4379 59814
rect 4435 59812 4459 59814
rect 4515 59812 4521 59814
rect 4213 59792 4521 59812
rect 4213 58780 4521 58800
rect 4213 58778 4219 58780
rect 4275 58778 4299 58780
rect 4355 58778 4379 58780
rect 4435 58778 4459 58780
rect 4515 58778 4521 58780
rect 4275 58726 4277 58778
rect 4457 58726 4459 58778
rect 4213 58724 4219 58726
rect 4275 58724 4299 58726
rect 4355 58724 4379 58726
rect 4435 58724 4459 58726
rect 4515 58724 4521 58726
rect 4213 58704 4521 58724
rect 4068 58064 4120 58070
rect 4068 58006 4120 58012
rect 4068 57928 4120 57934
rect 4068 57870 4120 57876
rect 4080 56846 4108 57870
rect 4213 57692 4521 57712
rect 4213 57690 4219 57692
rect 4275 57690 4299 57692
rect 4355 57690 4379 57692
rect 4435 57690 4459 57692
rect 4515 57690 4521 57692
rect 4275 57638 4277 57690
rect 4457 57638 4459 57690
rect 4213 57636 4219 57638
rect 4275 57636 4299 57638
rect 4355 57636 4379 57638
rect 4435 57636 4459 57638
rect 4515 57636 4521 57638
rect 4213 57616 4521 57636
rect 4068 56840 4120 56846
rect 4068 56782 4120 56788
rect 4213 56604 4521 56624
rect 4213 56602 4219 56604
rect 4275 56602 4299 56604
rect 4355 56602 4379 56604
rect 4435 56602 4459 56604
rect 4515 56602 4521 56604
rect 4275 56550 4277 56602
rect 4457 56550 4459 56602
rect 4213 56548 4219 56550
rect 4275 56548 4299 56550
rect 4355 56548 4379 56550
rect 4435 56548 4459 56550
rect 4515 56548 4521 56550
rect 4213 56528 4521 56548
rect 4213 55516 4521 55536
rect 4213 55514 4219 55516
rect 4275 55514 4299 55516
rect 4355 55514 4379 55516
rect 4435 55514 4459 55516
rect 4515 55514 4521 55516
rect 4275 55462 4277 55514
rect 4457 55462 4459 55514
rect 4213 55460 4219 55462
rect 4275 55460 4299 55462
rect 4355 55460 4379 55462
rect 4435 55460 4459 55462
rect 4515 55460 4521 55462
rect 4213 55440 4521 55460
rect 4213 54428 4521 54448
rect 4213 54426 4219 54428
rect 4275 54426 4299 54428
rect 4355 54426 4379 54428
rect 4435 54426 4459 54428
rect 4515 54426 4521 54428
rect 4275 54374 4277 54426
rect 4457 54374 4459 54426
rect 4213 54372 4219 54374
rect 4275 54372 4299 54374
rect 4355 54372 4379 54374
rect 4435 54372 4459 54374
rect 4515 54372 4521 54374
rect 4213 54352 4521 54372
rect 4213 53340 4521 53360
rect 4213 53338 4219 53340
rect 4275 53338 4299 53340
rect 4355 53338 4379 53340
rect 4435 53338 4459 53340
rect 4515 53338 4521 53340
rect 4275 53286 4277 53338
rect 4457 53286 4459 53338
rect 4213 53284 4219 53286
rect 4275 53284 4299 53286
rect 4355 53284 4379 53286
rect 4435 53284 4459 53286
rect 4515 53284 4521 53286
rect 4213 53264 4521 53284
rect 4213 52252 4521 52272
rect 4213 52250 4219 52252
rect 4275 52250 4299 52252
rect 4355 52250 4379 52252
rect 4435 52250 4459 52252
rect 4515 52250 4521 52252
rect 4275 52198 4277 52250
rect 4457 52198 4459 52250
rect 4213 52196 4219 52198
rect 4275 52196 4299 52198
rect 4355 52196 4379 52198
rect 4435 52196 4459 52198
rect 4515 52196 4521 52198
rect 4213 52176 4521 52196
rect 4213 51164 4521 51184
rect 4213 51162 4219 51164
rect 4275 51162 4299 51164
rect 4355 51162 4379 51164
rect 4435 51162 4459 51164
rect 4515 51162 4521 51164
rect 4275 51110 4277 51162
rect 4457 51110 4459 51162
rect 4213 51108 4219 51110
rect 4275 51108 4299 51110
rect 4355 51108 4379 51110
rect 4435 51108 4459 51110
rect 4515 51108 4521 51110
rect 4213 51088 4521 51108
rect 4160 50924 4212 50930
rect 4160 50866 4212 50872
rect 4172 50250 4200 50866
rect 4632 50425 4660 63854
rect 4988 59560 5040 59566
rect 4988 59502 5040 59508
rect 4896 57520 4948 57526
rect 4896 57462 4948 57468
rect 4804 55888 4856 55894
rect 4804 55830 4856 55836
rect 4712 54664 4764 54670
rect 4712 54606 4764 54612
rect 4618 50416 4674 50425
rect 4618 50351 4674 50360
rect 4160 50244 4212 50250
rect 4160 50186 4212 50192
rect 4620 50244 4672 50250
rect 4620 50186 4672 50192
rect 4213 50076 4521 50096
rect 4213 50074 4219 50076
rect 4275 50074 4299 50076
rect 4355 50074 4379 50076
rect 4435 50074 4459 50076
rect 4515 50074 4521 50076
rect 4275 50022 4277 50074
rect 4457 50022 4459 50074
rect 4213 50020 4219 50022
rect 4275 50020 4299 50022
rect 4355 50020 4379 50022
rect 4435 50020 4459 50022
rect 4515 50020 4521 50022
rect 4213 50000 4521 50020
rect 3988 49830 4108 49858
rect 3976 49768 4028 49774
rect 3976 49710 4028 49716
rect 3884 43444 3936 43450
rect 3884 43386 3936 43392
rect 3884 43308 3936 43314
rect 3884 43250 3936 43256
rect 3700 42696 3752 42702
rect 3700 42638 3752 42644
rect 3792 41744 3844 41750
rect 3792 41686 3844 41692
rect 3608 41540 3660 41546
rect 3608 41482 3660 41488
rect 3606 41440 3662 41449
rect 3606 41375 3662 41384
rect 3516 39092 3568 39098
rect 3516 39034 3568 39040
rect 3620 39030 3648 41375
rect 3608 39024 3660 39030
rect 3608 38966 3660 38972
rect 3516 38888 3568 38894
rect 3516 38830 3568 38836
rect 3424 38752 3476 38758
rect 3424 38694 3476 38700
rect 3436 38457 3464 38694
rect 3422 38448 3478 38457
rect 3422 38383 3478 38392
rect 3424 38208 3476 38214
rect 3424 38150 3476 38156
rect 3436 37874 3464 38150
rect 3424 37868 3476 37874
rect 3424 37810 3476 37816
rect 3160 34326 3372 34354
rect 3056 33856 3108 33862
rect 3056 33798 3108 33804
rect 2964 32904 3016 32910
rect 2964 32846 3016 32852
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 2780 31952 2832 31958
rect 2780 31894 2832 31900
rect 2504 31816 2556 31822
rect 2504 31758 2556 31764
rect 2504 31680 2556 31686
rect 2504 31622 2556 31628
rect 2412 31136 2464 31142
rect 2412 31078 2464 31084
rect 2320 28756 2372 28762
rect 2320 28698 2372 28704
rect 2424 28234 2452 31078
rect 2516 28694 2544 31622
rect 2792 31521 2820 31894
rect 2778 31512 2834 31521
rect 2778 31447 2834 31456
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2976 30818 3004 32846
rect 3160 31686 3188 34326
rect 3436 34218 3464 37810
rect 3344 34190 3464 34218
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 3252 32910 3280 33934
rect 3344 33386 3372 34190
rect 3528 33658 3556 38830
rect 3700 38752 3752 38758
rect 3700 38694 3752 38700
rect 3608 38344 3660 38350
rect 3606 38312 3608 38321
rect 3660 38312 3662 38321
rect 3606 38247 3662 38256
rect 3620 37806 3648 38247
rect 3608 37800 3660 37806
rect 3608 37742 3660 37748
rect 3608 36100 3660 36106
rect 3608 36042 3660 36048
rect 3620 35170 3648 36042
rect 3712 35698 3740 38694
rect 3700 35692 3752 35698
rect 3700 35634 3752 35640
rect 3620 35142 3740 35170
rect 3608 35080 3660 35086
rect 3608 35022 3660 35028
rect 3516 33652 3568 33658
rect 3516 33594 3568 33600
rect 3514 33552 3570 33561
rect 3424 33516 3476 33522
rect 3514 33487 3570 33496
rect 3424 33458 3476 33464
rect 3332 33380 3384 33386
rect 3332 33322 3384 33328
rect 3240 32904 3292 32910
rect 3240 32846 3292 32852
rect 3252 32434 3280 32846
rect 3240 32428 3292 32434
rect 3240 32370 3292 32376
rect 3148 31680 3200 31686
rect 3148 31622 3200 31628
rect 3056 31340 3108 31346
rect 3056 31282 3108 31288
rect 3068 30920 3096 31282
rect 3068 30892 3188 30920
rect 2596 30796 2648 30802
rect 2976 30790 3096 30818
rect 2596 30738 2648 30744
rect 2608 30326 2636 30738
rect 2964 30660 3016 30666
rect 2964 30602 3016 30608
rect 2596 30320 2648 30326
rect 2596 30262 2648 30268
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 2976 29306 3004 30602
rect 3068 30274 3096 30790
rect 3160 30394 3188 30892
rect 3148 30388 3200 30394
rect 3148 30330 3200 30336
rect 3068 30246 3188 30274
rect 3056 30048 3108 30054
rect 3056 29990 3108 29996
rect 2964 29300 3016 29306
rect 2964 29242 3016 29248
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 3068 28762 3096 29990
rect 3160 28801 3188 30246
rect 3252 29646 3280 32370
rect 3436 31754 3464 33458
rect 3344 31726 3464 31754
rect 3240 29640 3292 29646
rect 3240 29582 3292 29588
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 3146 28792 3202 28801
rect 3056 28756 3108 28762
rect 3146 28727 3202 28736
rect 3056 28698 3108 28704
rect 2504 28688 2556 28694
rect 3252 28665 3280 29106
rect 2504 28630 2556 28636
rect 3238 28656 3294 28665
rect 3238 28591 3294 28600
rect 2872 28552 2924 28558
rect 2870 28520 2872 28529
rect 2924 28520 2926 28529
rect 2870 28455 2926 28464
rect 3240 28484 3292 28490
rect 3240 28426 3292 28432
rect 2424 28206 2544 28234
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2424 27713 2452 28018
rect 2410 27704 2466 27713
rect 2410 27639 2466 27648
rect 2240 27526 2452 27554
rect 2148 27390 2360 27418
rect 2136 27328 2188 27334
rect 2136 27270 2188 27276
rect 2148 25786 2176 27270
rect 2228 26376 2280 26382
rect 2228 26318 2280 26324
rect 2240 26042 2268 26318
rect 2228 26036 2280 26042
rect 2228 25978 2280 25984
rect 2148 25758 2268 25786
rect 2136 25696 2188 25702
rect 2136 25638 2188 25644
rect 2148 24818 2176 25638
rect 2136 24812 2188 24818
rect 2136 24754 2188 24760
rect 2240 22778 2268 25758
rect 2332 24138 2360 27390
rect 2320 24132 2372 24138
rect 2320 24074 2372 24080
rect 2424 23798 2452 27526
rect 2516 27334 2544 28206
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2976 27606 3004 27950
rect 2964 27600 3016 27606
rect 2964 27542 3016 27548
rect 2964 27464 3016 27470
rect 2964 27406 3016 27412
rect 2504 27328 2556 27334
rect 2976 27305 3004 27406
rect 2504 27270 2556 27276
rect 2962 27296 3018 27305
rect 2962 27231 3018 27240
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 3148 26988 3200 26994
rect 3148 26930 3200 26936
rect 2516 26586 2544 26930
rect 3160 26897 3188 26930
rect 3146 26888 3202 26897
rect 3146 26823 3202 26832
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 2504 26580 2556 26586
rect 2504 26522 2556 26528
rect 2688 26444 2740 26450
rect 2688 26386 2740 26392
rect 2700 26042 2728 26386
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 2688 26036 2740 26042
rect 2688 25978 2740 25984
rect 3068 25945 3096 26318
rect 3054 25936 3110 25945
rect 2872 25900 2924 25906
rect 3054 25871 3110 25880
rect 2872 25842 2924 25848
rect 2884 25809 2912 25842
rect 2870 25800 2926 25809
rect 2870 25735 2926 25744
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2780 25288 2832 25294
rect 2780 25230 2832 25236
rect 2792 24721 2820 25230
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2778 24712 2834 24721
rect 2778 24647 2834 24656
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2504 24132 2556 24138
rect 2504 24074 2556 24080
rect 2412 23792 2464 23798
rect 2412 23734 2464 23740
rect 2424 23118 2452 23734
rect 2516 23730 2544 24074
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2424 22658 2452 23054
rect 2516 22778 2544 23666
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2872 23248 2924 23254
rect 2976 23225 3004 24754
rect 3252 24682 3280 28426
rect 3344 26432 3372 31726
rect 3424 31272 3476 31278
rect 3424 31214 3476 31220
rect 3436 29850 3464 31214
rect 3528 30938 3556 33487
rect 3516 30932 3568 30938
rect 3516 30874 3568 30880
rect 3516 30728 3568 30734
rect 3516 30670 3568 30676
rect 3424 29844 3476 29850
rect 3424 29786 3476 29792
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3436 27538 3464 29582
rect 3424 27532 3476 27538
rect 3424 27474 3476 27480
rect 3344 26404 3464 26432
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 3240 24676 3292 24682
rect 3240 24618 3292 24624
rect 3240 24064 3292 24070
rect 3240 24006 3292 24012
rect 3252 23730 3280 24006
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 2872 23190 2924 23196
rect 2962 23216 3018 23225
rect 2688 23180 2740 23186
rect 2688 23122 2740 23128
rect 2504 22772 2556 22778
rect 2504 22714 2556 22720
rect 2136 22636 2188 22642
rect 2136 22578 2188 22584
rect 2332 22630 2544 22658
rect 2148 18834 2176 22578
rect 2332 22030 2360 22630
rect 2516 22574 2544 22630
rect 2504 22568 2556 22574
rect 2504 22510 2556 22516
rect 2700 22506 2728 23122
rect 2884 22710 2912 23190
rect 2962 23151 3018 23160
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2412 22500 2464 22506
rect 2412 22442 2464 22448
rect 2688 22500 2740 22506
rect 2688 22442 2740 22448
rect 2424 22030 2452 22442
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2228 21412 2280 21418
rect 2228 21354 2280 21360
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 2240 18358 2268 21354
rect 2424 20210 2452 21966
rect 2976 21690 3004 23054
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 3068 22234 3096 22714
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 3160 21729 3188 21966
rect 3146 21720 3202 21729
rect 2964 21684 3016 21690
rect 3146 21655 3202 21664
rect 2964 21626 3016 21632
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2516 20942 2544 21286
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2792 20369 2820 20402
rect 2964 20392 3016 20398
rect 2778 20360 2834 20369
rect 2964 20334 3016 20340
rect 2778 20295 2834 20304
rect 2332 20182 2452 20210
rect 2228 18352 2280 18358
rect 1964 17190 2084 17218
rect 2148 18312 2228 18340
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13569 1716 14350
rect 1872 14056 1900 14962
rect 1780 14028 1900 14056
rect 1674 13560 1730 13569
rect 1674 13495 1730 13504
rect 1780 13258 1808 14028
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 13252 1820 13258
rect 1768 13194 1820 13200
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1504 12406 1624 12434
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1306 11792 1362 11801
rect 1306 11727 1362 11736
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 10985 1348 11630
rect 1412 11393 1440 12174
rect 1398 11384 1454 11393
rect 1398 11319 1454 11328
rect 1504 11218 1532 12406
rect 1780 11762 1808 12922
rect 1872 12617 1900 13874
rect 1858 12608 1914 12617
rect 1858 12543 1914 12552
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1320 10033 1348 10542
rect 1412 10441 1440 11086
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1400 10056 1452 10062
rect 1306 10024 1362 10033
rect 1400 9998 1452 10004
rect 1306 9959 1362 9968
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9217 1440 9454
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1584 8900 1636 8906
rect 1584 8842 1636 8848
rect 1596 8634 1624 8842
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1216 7472 1268 7478
rect 1412 7449 1440 7822
rect 1216 7414 1268 7420
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1504 6798 1532 8434
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1412 6633 1440 6734
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 1320 3641 1348 5646
rect 1412 4865 1440 6258
rect 1504 5914 1532 6734
rect 1596 6458 1624 8434
rect 1872 7886 1900 8910
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1596 5234 1624 5646
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 1306 3632 1362 3641
rect 1306 3567 1362 3576
rect 1398 3224 1454 3233
rect 1398 3159 1454 3168
rect 1412 2446 1440 3159
rect 1596 2650 1624 5170
rect 1964 4214 1992 17190
rect 2148 16250 2176 18312
rect 2228 18294 2280 18300
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 16658 2268 16934
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2332 16522 2360 20182
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 2976 19961 3004 20334
rect 2962 19952 3018 19961
rect 2962 19887 3018 19896
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2792 19281 2820 19790
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 2778 19272 2834 19281
rect 2778 19207 2834 19216
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2424 18426 2452 18702
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2412 18284 2464 18290
rect 2412 18226 2464 18232
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2424 16266 2452 18226
rect 2516 17678 2544 19110
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2700 18290 2728 18702
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2976 18193 3004 19314
rect 3068 18358 3096 21490
rect 3148 20868 3200 20874
rect 3148 20810 3200 20816
rect 3160 20602 3188 20810
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3160 19553 3188 19790
rect 3146 19544 3202 19553
rect 3146 19479 3202 19488
rect 3252 19394 3280 22986
rect 3160 19366 3280 19394
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 2962 18184 3018 18193
rect 2962 18119 3018 18128
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 17105 2912 17138
rect 2870 17096 2926 17105
rect 2870 17031 2926 17040
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2240 16238 2452 16266
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2056 15706 2084 15982
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2056 13394 2084 15642
rect 2240 15586 2268 16238
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2148 15558 2268 15586
rect 2148 15162 2176 15558
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2136 14884 2188 14890
rect 2136 14826 2188 14832
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 2056 12306 2084 13194
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2148 10674 2176 14826
rect 2240 14793 2268 15438
rect 2226 14784 2282 14793
rect 2226 14719 2282 14728
rect 2332 14634 2360 16050
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 14958 2452 15846
rect 2516 15434 2544 16458
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2608 15978 2636 16390
rect 2792 16017 2820 16526
rect 2778 16008 2834 16017
rect 2596 15972 2648 15978
rect 2778 15943 2834 15952
rect 2596 15914 2648 15920
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2884 15201 2912 15438
rect 2870 15192 2926 15201
rect 3068 15162 3096 18294
rect 3160 16574 3188 19366
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3252 17746 3280 18022
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3160 16546 3280 16574
rect 3252 16046 3280 16546
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 2870 15127 2926 15136
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2412 14952 2464 14958
rect 2412 14894 2464 14900
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2240 14606 2360 14634
rect 2240 12850 2268 14606
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2240 11150 2268 11698
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 8498 2176 9998
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2056 7041 2084 7346
rect 2042 7032 2098 7041
rect 2042 6967 2098 6976
rect 2240 6458 2268 11086
rect 2332 9586 2360 13942
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2424 9042 2452 9522
rect 2516 9450 2544 14758
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 2976 14074 3004 14962
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3160 13977 3188 14350
rect 3146 13968 3202 13977
rect 3146 13903 3202 13912
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 13025 2820 13194
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 7954 2452 8978
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8498 2912 8910
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5273 2084 6258
rect 2042 5264 2098 5273
rect 2042 5199 2098 5208
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 3194 2268 3470
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2332 2650 2360 5170
rect 2516 3738 2544 7822
rect 2792 7546 2820 7958
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2976 6914 3004 10474
rect 3068 9058 3096 10610
rect 3160 10130 3188 13806
rect 3252 13462 3280 15982
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3344 13002 3372 26250
rect 3436 24614 3464 26404
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3424 24268 3476 24274
rect 3424 24210 3476 24216
rect 3436 23662 3464 24210
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3436 23254 3464 23598
rect 3424 23248 3476 23254
rect 3424 23190 3476 23196
rect 3436 22778 3464 23190
rect 3528 22778 3556 30670
rect 3424 22772 3476 22778
rect 3424 22714 3476 22720
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3436 22545 3464 22578
rect 3620 22556 3648 35022
rect 3712 32910 3740 35142
rect 3700 32904 3752 32910
rect 3700 32846 3752 32852
rect 3700 32768 3752 32774
rect 3700 32710 3752 32716
rect 3712 25498 3740 32710
rect 3804 32065 3832 41686
rect 3896 32774 3924 43250
rect 3988 41449 4016 49710
rect 4080 46102 4108 49830
rect 4632 49638 4660 50186
rect 4620 49632 4672 49638
rect 4620 49574 4672 49580
rect 4620 49224 4672 49230
rect 4620 49166 4672 49172
rect 4213 48988 4521 49008
rect 4213 48986 4219 48988
rect 4275 48986 4299 48988
rect 4355 48986 4379 48988
rect 4435 48986 4459 48988
rect 4515 48986 4521 48988
rect 4275 48934 4277 48986
rect 4457 48934 4459 48986
rect 4213 48932 4219 48934
rect 4275 48932 4299 48934
rect 4355 48932 4379 48934
rect 4435 48932 4459 48934
rect 4515 48932 4521 48934
rect 4213 48912 4521 48932
rect 4526 48784 4582 48793
rect 4526 48719 4582 48728
rect 4540 48210 4568 48719
rect 4528 48204 4580 48210
rect 4528 48146 4580 48152
rect 4213 47900 4521 47920
rect 4213 47898 4219 47900
rect 4275 47898 4299 47900
rect 4355 47898 4379 47900
rect 4435 47898 4459 47900
rect 4515 47898 4521 47900
rect 4275 47846 4277 47898
rect 4457 47846 4459 47898
rect 4213 47844 4219 47846
rect 4275 47844 4299 47846
rect 4355 47844 4379 47846
rect 4435 47844 4459 47846
rect 4515 47844 4521 47846
rect 4213 47824 4521 47844
rect 4213 46812 4521 46832
rect 4213 46810 4219 46812
rect 4275 46810 4299 46812
rect 4355 46810 4379 46812
rect 4435 46810 4459 46812
rect 4515 46810 4521 46812
rect 4275 46758 4277 46810
rect 4457 46758 4459 46810
rect 4213 46756 4219 46758
rect 4275 46756 4299 46758
rect 4355 46756 4379 46758
rect 4435 46756 4459 46758
rect 4515 46756 4521 46758
rect 4213 46736 4521 46756
rect 4632 46594 4660 49166
rect 4448 46566 4660 46594
rect 4068 46096 4120 46102
rect 4448 46073 4476 46566
rect 4724 46458 4752 54606
rect 4540 46430 4752 46458
rect 4540 46102 4568 46430
rect 4620 46368 4672 46374
rect 4816 46322 4844 55830
rect 4620 46310 4672 46316
rect 4528 46096 4580 46102
rect 4068 46038 4120 46044
rect 4434 46064 4490 46073
rect 4528 46038 4580 46044
rect 4434 45999 4490 46008
rect 4213 45724 4521 45744
rect 4213 45722 4219 45724
rect 4275 45722 4299 45724
rect 4355 45722 4379 45724
rect 4435 45722 4459 45724
rect 4515 45722 4521 45724
rect 4275 45670 4277 45722
rect 4457 45670 4459 45722
rect 4213 45668 4219 45670
rect 4275 45668 4299 45670
rect 4355 45668 4379 45670
rect 4435 45668 4459 45670
rect 4515 45668 4521 45670
rect 4213 45648 4521 45668
rect 4068 45076 4120 45082
rect 4068 45018 4120 45024
rect 3974 41440 4030 41449
rect 3974 41375 4030 41384
rect 3976 41268 4028 41274
rect 3976 41210 4028 41216
rect 3988 36258 4016 41210
rect 4080 41138 4108 45018
rect 4213 44636 4521 44656
rect 4213 44634 4219 44636
rect 4275 44634 4299 44636
rect 4355 44634 4379 44636
rect 4435 44634 4459 44636
rect 4515 44634 4521 44636
rect 4275 44582 4277 44634
rect 4457 44582 4459 44634
rect 4213 44580 4219 44582
rect 4275 44580 4299 44582
rect 4355 44580 4379 44582
rect 4435 44580 4459 44582
rect 4515 44580 4521 44582
rect 4213 44560 4521 44580
rect 4158 44432 4214 44441
rect 4158 44367 4160 44376
rect 4212 44367 4214 44376
rect 4160 44338 4212 44344
rect 4172 43790 4200 44338
rect 4160 43784 4212 43790
rect 4160 43726 4212 43732
rect 4213 43548 4521 43568
rect 4213 43546 4219 43548
rect 4275 43546 4299 43548
rect 4355 43546 4379 43548
rect 4435 43546 4459 43548
rect 4515 43546 4521 43548
rect 4275 43494 4277 43546
rect 4457 43494 4459 43546
rect 4213 43492 4219 43494
rect 4275 43492 4299 43494
rect 4355 43492 4379 43494
rect 4435 43492 4459 43494
rect 4515 43492 4521 43494
rect 4213 43472 4521 43492
rect 4160 43308 4212 43314
rect 4160 43250 4212 43256
rect 4172 43110 4200 43250
rect 4160 43104 4212 43110
rect 4160 43046 4212 43052
rect 4172 42906 4200 43046
rect 4160 42900 4212 42906
rect 4160 42842 4212 42848
rect 4213 42460 4521 42480
rect 4213 42458 4219 42460
rect 4275 42458 4299 42460
rect 4355 42458 4379 42460
rect 4435 42458 4459 42460
rect 4515 42458 4521 42460
rect 4275 42406 4277 42458
rect 4457 42406 4459 42458
rect 4213 42404 4219 42406
rect 4275 42404 4299 42406
rect 4355 42404 4379 42406
rect 4435 42404 4459 42406
rect 4515 42404 4521 42406
rect 4213 42384 4521 42404
rect 4213 41372 4521 41392
rect 4213 41370 4219 41372
rect 4275 41370 4299 41372
rect 4355 41370 4379 41372
rect 4435 41370 4459 41372
rect 4515 41370 4521 41372
rect 4275 41318 4277 41370
rect 4457 41318 4459 41370
rect 4213 41316 4219 41318
rect 4275 41316 4299 41318
rect 4355 41316 4379 41318
rect 4435 41316 4459 41318
rect 4515 41316 4521 41318
rect 4213 41296 4521 41316
rect 4068 41132 4120 41138
rect 4068 41074 4120 41080
rect 4213 40284 4521 40304
rect 4213 40282 4219 40284
rect 4275 40282 4299 40284
rect 4355 40282 4379 40284
rect 4435 40282 4459 40284
rect 4515 40282 4521 40284
rect 4275 40230 4277 40282
rect 4457 40230 4459 40282
rect 4213 40228 4219 40230
rect 4275 40228 4299 40230
rect 4355 40228 4379 40230
rect 4435 40228 4459 40230
rect 4515 40228 4521 40230
rect 4213 40208 4521 40228
rect 4213 39196 4521 39216
rect 4213 39194 4219 39196
rect 4275 39194 4299 39196
rect 4355 39194 4379 39196
rect 4435 39194 4459 39196
rect 4515 39194 4521 39196
rect 4275 39142 4277 39194
rect 4457 39142 4459 39194
rect 4213 39140 4219 39142
rect 4275 39140 4299 39142
rect 4355 39140 4379 39142
rect 4435 39140 4459 39142
rect 4515 39140 4521 39142
rect 4213 39120 4521 39140
rect 4068 38956 4120 38962
rect 4068 38898 4120 38904
rect 4080 38350 4108 38898
rect 4068 38344 4120 38350
rect 4068 38286 4120 38292
rect 4213 38108 4521 38128
rect 4213 38106 4219 38108
rect 4275 38106 4299 38108
rect 4355 38106 4379 38108
rect 4435 38106 4459 38108
rect 4515 38106 4521 38108
rect 4275 38054 4277 38106
rect 4457 38054 4459 38106
rect 4213 38052 4219 38054
rect 4275 38052 4299 38054
rect 4355 38052 4379 38054
rect 4435 38052 4459 38054
rect 4515 38052 4521 38054
rect 4213 38032 4521 38052
rect 4632 37194 4660 46310
rect 4724 46294 4844 46322
rect 4724 46034 4752 46294
rect 4804 46164 4856 46170
rect 4804 46106 4856 46112
rect 4712 46028 4764 46034
rect 4712 45970 4764 45976
rect 4712 45892 4764 45898
rect 4712 45834 4764 45840
rect 4620 37188 4672 37194
rect 4620 37130 4672 37136
rect 4213 37020 4521 37040
rect 4213 37018 4219 37020
rect 4275 37018 4299 37020
rect 4355 37018 4379 37020
rect 4435 37018 4459 37020
rect 4515 37018 4521 37020
rect 4275 36966 4277 37018
rect 4457 36966 4459 37018
rect 4213 36964 4219 36966
rect 4275 36964 4299 36966
rect 4355 36964 4379 36966
rect 4435 36964 4459 36966
rect 4515 36964 4521 36966
rect 4213 36944 4521 36964
rect 3988 36230 4108 36258
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3988 35086 4016 36110
rect 3976 35080 4028 35086
rect 3976 35022 4028 35028
rect 3988 33998 4016 35022
rect 3976 33992 4028 33998
rect 3976 33934 4028 33940
rect 4080 32994 4108 36230
rect 4213 35932 4521 35952
rect 4213 35930 4219 35932
rect 4275 35930 4299 35932
rect 4355 35930 4379 35932
rect 4435 35930 4459 35932
rect 4515 35930 4521 35932
rect 4275 35878 4277 35930
rect 4457 35878 4459 35930
rect 4213 35876 4219 35878
rect 4275 35876 4299 35878
rect 4355 35876 4379 35878
rect 4435 35876 4459 35878
rect 4515 35876 4521 35878
rect 4213 35856 4521 35876
rect 4724 35834 4752 45834
rect 4816 40118 4844 46106
rect 4804 40112 4856 40118
rect 4804 40054 4856 40060
rect 4908 38010 4936 57462
rect 5000 46170 5028 59502
rect 4988 46164 5040 46170
rect 4988 46106 5040 46112
rect 4988 46028 5040 46034
rect 4988 45970 5040 45976
rect 4896 38004 4948 38010
rect 4896 37946 4948 37952
rect 5000 36310 5028 45970
rect 5092 45082 5120 71062
rect 5172 68128 5224 68134
rect 5172 68070 5224 68076
rect 5184 49774 5212 68070
rect 5356 57248 5408 57254
rect 5356 57190 5408 57196
rect 5264 56296 5316 56302
rect 5264 56238 5316 56244
rect 5172 49768 5224 49774
rect 5172 49710 5224 49716
rect 5172 49632 5224 49638
rect 5172 49574 5224 49580
rect 5184 45626 5212 49574
rect 5172 45620 5224 45626
rect 5172 45562 5224 45568
rect 5170 45520 5226 45529
rect 5170 45455 5226 45464
rect 5080 45076 5132 45082
rect 5080 45018 5132 45024
rect 5078 42528 5134 42537
rect 5078 42463 5134 42472
rect 4988 36304 5040 36310
rect 4988 36246 5040 36252
rect 4712 35828 4764 35834
rect 4712 35770 4764 35776
rect 4213 34844 4521 34864
rect 4213 34842 4219 34844
rect 4275 34842 4299 34844
rect 4355 34842 4379 34844
rect 4435 34842 4459 34844
rect 4515 34842 4521 34844
rect 4275 34790 4277 34842
rect 4457 34790 4459 34842
rect 4213 34788 4219 34790
rect 4275 34788 4299 34790
rect 4355 34788 4379 34790
rect 4435 34788 4459 34790
rect 4515 34788 4521 34790
rect 4213 34768 4521 34788
rect 4620 33924 4672 33930
rect 4620 33866 4672 33872
rect 4213 33756 4521 33776
rect 4213 33754 4219 33756
rect 4275 33754 4299 33756
rect 4355 33754 4379 33756
rect 4435 33754 4459 33756
rect 4515 33754 4521 33756
rect 4275 33702 4277 33754
rect 4457 33702 4459 33754
rect 4213 33700 4219 33702
rect 4275 33700 4299 33702
rect 4355 33700 4379 33702
rect 4435 33700 4459 33702
rect 4515 33700 4521 33702
rect 4213 33680 4521 33700
rect 3988 32966 4108 32994
rect 3884 32768 3936 32774
rect 3884 32710 3936 32716
rect 3988 32502 4016 32966
rect 4068 32836 4120 32842
rect 4068 32778 4120 32784
rect 3976 32496 4028 32502
rect 3976 32438 4028 32444
rect 3790 32056 3846 32065
rect 3790 31991 3846 32000
rect 3792 31884 3844 31890
rect 3792 31826 3844 31832
rect 3804 30938 3832 31826
rect 3792 30932 3844 30938
rect 3792 30874 3844 30880
rect 3976 30728 4028 30734
rect 3976 30670 4028 30676
rect 3988 30297 4016 30670
rect 3974 30288 4030 30297
rect 3974 30223 4030 30232
rect 3790 30152 3846 30161
rect 3790 30087 3846 30096
rect 3884 30116 3936 30122
rect 3700 25492 3752 25498
rect 3700 25434 3752 25440
rect 3700 24064 3752 24070
rect 3700 24006 3752 24012
rect 3422 22536 3478 22545
rect 3422 22471 3478 22480
rect 3528 22528 3648 22556
rect 3528 22386 3556 22528
rect 3712 22488 3740 24006
rect 3436 22358 3556 22386
rect 3620 22460 3740 22488
rect 3436 20330 3464 22358
rect 3620 22094 3648 22460
rect 3804 22386 3832 30087
rect 3884 30058 3936 30064
rect 3896 29753 3924 30058
rect 3882 29744 3938 29753
rect 3882 29679 3938 29688
rect 3976 29640 4028 29646
rect 3976 29582 4028 29588
rect 3884 29504 3936 29510
rect 3884 29446 3936 29452
rect 3896 23610 3924 29446
rect 3988 29345 4016 29582
rect 3974 29336 4030 29345
rect 3974 29271 4030 29280
rect 3976 27532 4028 27538
rect 3976 27474 4028 27480
rect 3988 24342 4016 27474
rect 3976 24336 4028 24342
rect 3976 24278 4028 24284
rect 3976 24200 4028 24206
rect 3976 24142 4028 24148
rect 3988 23769 4016 24142
rect 3974 23760 4030 23769
rect 3974 23695 4030 23704
rect 3896 23582 4016 23610
rect 3884 23316 3936 23322
rect 3884 23258 3936 23264
rect 3528 22066 3648 22094
rect 3712 22358 3832 22386
rect 3424 20324 3476 20330
rect 3424 20266 3476 20272
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3436 17785 3464 18226
rect 3422 17776 3478 17785
rect 3422 17711 3478 17720
rect 3252 12974 3372 13002
rect 3252 11830 3280 12974
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3436 11762 3464 12786
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3148 10124 3200 10130
rect 3148 10066 3200 10072
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3252 9178 3280 9522
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3068 9030 3280 9058
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3068 8809 3096 8910
rect 3054 8800 3110 8809
rect 3054 8735 3110 8744
rect 3160 7954 3188 8910
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3252 6914 3280 9030
rect 3436 8242 3464 11698
rect 3528 8974 3556 22066
rect 3606 21992 3662 22001
rect 3606 21927 3662 21936
rect 3620 19242 3648 21927
rect 3712 21146 3740 22358
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3804 21026 3832 22170
rect 3712 20998 3832 21026
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3620 11354 3648 11494
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 10282 3740 20998
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 3804 20058 3832 20810
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3804 17882 3832 18158
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 3896 16574 3924 23258
rect 3988 21026 4016 23582
rect 4080 21146 4108 32778
rect 4213 32668 4521 32688
rect 4213 32666 4219 32668
rect 4275 32666 4299 32668
rect 4355 32666 4379 32668
rect 4435 32666 4459 32668
rect 4515 32666 4521 32668
rect 4275 32614 4277 32666
rect 4457 32614 4459 32666
rect 4213 32612 4219 32614
rect 4275 32612 4299 32614
rect 4355 32612 4379 32614
rect 4435 32612 4459 32614
rect 4515 32612 4521 32614
rect 4213 32592 4521 32612
rect 4213 31580 4521 31600
rect 4213 31578 4219 31580
rect 4275 31578 4299 31580
rect 4355 31578 4379 31580
rect 4435 31578 4459 31580
rect 4515 31578 4521 31580
rect 4275 31526 4277 31578
rect 4457 31526 4459 31578
rect 4213 31524 4219 31526
rect 4275 31524 4299 31526
rect 4355 31524 4379 31526
rect 4435 31524 4459 31526
rect 4515 31524 4521 31526
rect 4213 31504 4521 31524
rect 4213 30492 4521 30512
rect 4213 30490 4219 30492
rect 4275 30490 4299 30492
rect 4355 30490 4379 30492
rect 4435 30490 4459 30492
rect 4515 30490 4521 30492
rect 4275 30438 4277 30490
rect 4457 30438 4459 30490
rect 4213 30436 4219 30438
rect 4275 30436 4299 30438
rect 4355 30436 4379 30438
rect 4435 30436 4459 30438
rect 4515 30436 4521 30438
rect 4213 30416 4521 30436
rect 4632 29510 4660 33866
rect 4712 29572 4764 29578
rect 4712 29514 4764 29520
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4213 29404 4521 29424
rect 4213 29402 4219 29404
rect 4275 29402 4299 29404
rect 4355 29402 4379 29404
rect 4435 29402 4459 29404
rect 4515 29402 4521 29404
rect 4275 29350 4277 29402
rect 4457 29350 4459 29402
rect 4213 29348 4219 29350
rect 4275 29348 4299 29350
rect 4355 29348 4379 29350
rect 4435 29348 4459 29350
rect 4515 29348 4521 29350
rect 4213 29328 4521 29348
rect 4213 28316 4521 28336
rect 4213 28314 4219 28316
rect 4275 28314 4299 28316
rect 4355 28314 4379 28316
rect 4435 28314 4459 28316
rect 4515 28314 4521 28316
rect 4275 28262 4277 28314
rect 4457 28262 4459 28314
rect 4213 28260 4219 28262
rect 4275 28260 4299 28262
rect 4355 28260 4379 28262
rect 4435 28260 4459 28262
rect 4515 28260 4521 28262
rect 4213 28240 4521 28260
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4213 27228 4521 27248
rect 4213 27226 4219 27228
rect 4275 27226 4299 27228
rect 4355 27226 4379 27228
rect 4435 27226 4459 27228
rect 4515 27226 4521 27228
rect 4275 27174 4277 27226
rect 4457 27174 4459 27226
rect 4213 27172 4219 27174
rect 4275 27172 4299 27174
rect 4355 27172 4379 27174
rect 4435 27172 4459 27174
rect 4515 27172 4521 27174
rect 4213 27152 4521 27172
rect 4213 26140 4521 26160
rect 4213 26138 4219 26140
rect 4275 26138 4299 26140
rect 4355 26138 4379 26140
rect 4435 26138 4459 26140
rect 4515 26138 4521 26140
rect 4275 26086 4277 26138
rect 4457 26086 4459 26138
rect 4213 26084 4219 26086
rect 4275 26084 4299 26086
rect 4355 26084 4379 26086
rect 4435 26084 4459 26086
rect 4515 26084 4521 26086
rect 4213 26064 4521 26084
rect 4213 25052 4521 25072
rect 4213 25050 4219 25052
rect 4275 25050 4299 25052
rect 4355 25050 4379 25052
rect 4435 25050 4459 25052
rect 4515 25050 4521 25052
rect 4275 24998 4277 25050
rect 4457 24998 4459 25050
rect 4213 24996 4219 24998
rect 4275 24996 4299 24998
rect 4355 24996 4379 24998
rect 4435 24996 4459 24998
rect 4515 24996 4521 24998
rect 4213 24976 4521 24996
rect 4213 23964 4521 23984
rect 4213 23962 4219 23964
rect 4275 23962 4299 23964
rect 4355 23962 4379 23964
rect 4435 23962 4459 23964
rect 4515 23962 4521 23964
rect 4275 23910 4277 23962
rect 4457 23910 4459 23962
rect 4213 23908 4219 23910
rect 4275 23908 4299 23910
rect 4355 23908 4379 23910
rect 4435 23908 4459 23910
rect 4515 23908 4521 23910
rect 4213 23888 4521 23908
rect 4632 22982 4660 27406
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 4213 22876 4521 22896
rect 4213 22874 4219 22876
rect 4275 22874 4299 22876
rect 4355 22874 4379 22876
rect 4435 22874 4459 22876
rect 4515 22874 4521 22876
rect 4275 22822 4277 22874
rect 4457 22822 4459 22874
rect 4213 22820 4219 22822
rect 4275 22820 4299 22822
rect 4355 22820 4379 22822
rect 4435 22820 4459 22822
rect 4515 22820 4521 22822
rect 4213 22800 4521 22820
rect 4213 21788 4521 21808
rect 4213 21786 4219 21788
rect 4275 21786 4299 21788
rect 4355 21786 4379 21788
rect 4435 21786 4459 21788
rect 4515 21786 4521 21788
rect 4275 21734 4277 21786
rect 4457 21734 4459 21786
rect 4213 21732 4219 21734
rect 4275 21732 4299 21734
rect 4355 21732 4379 21734
rect 4435 21732 4459 21734
rect 4515 21732 4521 21734
rect 4213 21712 4521 21732
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 3988 20998 4108 21026
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3988 20777 4016 20878
rect 4080 20806 4108 20998
rect 4068 20800 4120 20806
rect 3974 20768 4030 20777
rect 4068 20742 4120 20748
rect 3974 20703 4030 20712
rect 4213 20700 4521 20720
rect 4213 20698 4219 20700
rect 4275 20698 4299 20700
rect 4355 20698 4379 20700
rect 4435 20698 4459 20700
rect 4515 20698 4521 20700
rect 4275 20646 4277 20698
rect 4457 20646 4459 20698
rect 4213 20644 4219 20646
rect 4275 20644 4299 20646
rect 4355 20644 4379 20646
rect 4435 20644 4459 20646
rect 4515 20644 4521 20646
rect 4213 20624 4521 20644
rect 4213 19612 4521 19632
rect 4213 19610 4219 19612
rect 4275 19610 4299 19612
rect 4355 19610 4379 19612
rect 4435 19610 4459 19612
rect 4515 19610 4521 19612
rect 4275 19558 4277 19610
rect 4457 19558 4459 19610
rect 4213 19556 4219 19558
rect 4275 19556 4299 19558
rect 4355 19556 4379 19558
rect 4435 19556 4459 19558
rect 4515 19556 4521 19558
rect 4213 19536 4521 19556
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3988 18601 4016 18702
rect 3974 18592 4030 18601
rect 3974 18527 4030 18536
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3988 17377 4016 17614
rect 3974 17368 4030 17377
rect 3974 17303 4030 17312
rect 3804 16546 3924 16574
rect 3804 12238 3832 16546
rect 3976 14408 4028 14414
rect 3974 14376 3976 14385
rect 4028 14376 4030 14385
rect 3974 14311 4030 14320
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3620 10254 3740 10282
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 8401 3556 8434
rect 3514 8392 3570 8401
rect 3514 8327 3570 8336
rect 3436 8214 3556 8242
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 2976 6886 3188 6914
rect 3252 6886 3372 6914
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2976 5817 3004 6258
rect 2962 5808 3018 5817
rect 2962 5743 3018 5752
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 2976 4690 3004 4966
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 3160 4010 3188 6886
rect 3344 6474 3372 6886
rect 3252 6446 3372 6474
rect 3252 5302 3280 6446
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 3344 6225 3372 6258
rect 3330 6216 3386 6225
rect 3330 6151 3386 6160
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3436 5234 3464 7890
rect 3528 6458 3556 8214
rect 3620 7410 3648 10254
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3712 8634 3740 9590
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 7698 3740 8366
rect 3804 8022 3832 12174
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3896 11150 3924 12106
rect 4080 11880 4108 18770
rect 4213 18524 4521 18544
rect 4213 18522 4219 18524
rect 4275 18522 4299 18524
rect 4355 18522 4379 18524
rect 4435 18522 4459 18524
rect 4515 18522 4521 18524
rect 4275 18470 4277 18522
rect 4457 18470 4459 18522
rect 4213 18468 4219 18470
rect 4275 18468 4299 18470
rect 4355 18468 4379 18470
rect 4435 18468 4459 18470
rect 4515 18468 4521 18470
rect 4213 18448 4521 18468
rect 4213 17436 4521 17456
rect 4213 17434 4219 17436
rect 4275 17434 4299 17436
rect 4355 17434 4379 17436
rect 4435 17434 4459 17436
rect 4515 17434 4521 17436
rect 4275 17382 4277 17434
rect 4457 17382 4459 17434
rect 4213 17380 4219 17382
rect 4275 17380 4299 17382
rect 4355 17380 4379 17382
rect 4435 17380 4459 17382
rect 4515 17380 4521 17382
rect 4213 17360 4521 17380
rect 4213 16348 4521 16368
rect 4213 16346 4219 16348
rect 4275 16346 4299 16348
rect 4355 16346 4379 16348
rect 4435 16346 4459 16348
rect 4515 16346 4521 16348
rect 4275 16294 4277 16346
rect 4457 16294 4459 16346
rect 4213 16292 4219 16294
rect 4275 16292 4299 16294
rect 4355 16292 4379 16294
rect 4435 16292 4459 16294
rect 4515 16292 4521 16294
rect 4213 16272 4521 16292
rect 4213 15260 4521 15280
rect 4213 15258 4219 15260
rect 4275 15258 4299 15260
rect 4355 15258 4379 15260
rect 4435 15258 4459 15260
rect 4515 15258 4521 15260
rect 4275 15206 4277 15258
rect 4457 15206 4459 15258
rect 4213 15204 4219 15206
rect 4275 15204 4299 15206
rect 4355 15204 4379 15206
rect 4435 15204 4459 15206
rect 4515 15204 4521 15206
rect 4213 15184 4521 15204
rect 4213 14172 4521 14192
rect 4213 14170 4219 14172
rect 4275 14170 4299 14172
rect 4355 14170 4379 14172
rect 4435 14170 4459 14172
rect 4515 14170 4521 14172
rect 4275 14118 4277 14170
rect 4457 14118 4459 14170
rect 4213 14116 4219 14118
rect 4275 14116 4299 14118
rect 4355 14116 4379 14118
rect 4435 14116 4459 14118
rect 4515 14116 4521 14118
rect 4213 14096 4521 14116
rect 4213 13084 4521 13104
rect 4213 13082 4219 13084
rect 4275 13082 4299 13084
rect 4355 13082 4379 13084
rect 4435 13082 4459 13084
rect 4515 13082 4521 13084
rect 4275 13030 4277 13082
rect 4457 13030 4459 13082
rect 4213 13028 4219 13030
rect 4275 13028 4299 13030
rect 4355 13028 4379 13030
rect 4435 13028 4459 13030
rect 4515 13028 4521 13030
rect 4213 13008 4521 13028
rect 4213 11996 4521 12016
rect 4213 11994 4219 11996
rect 4275 11994 4299 11996
rect 4355 11994 4379 11996
rect 4435 11994 4459 11996
rect 4515 11994 4521 11996
rect 4275 11942 4277 11994
rect 4457 11942 4459 11994
rect 4213 11940 4219 11942
rect 4275 11940 4299 11942
rect 4355 11940 4379 11942
rect 4435 11940 4459 11942
rect 4515 11940 4521 11942
rect 4213 11920 4521 11940
rect 3988 11852 4108 11880
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3792 7880 3844 7886
rect 3790 7848 3792 7857
rect 3844 7848 3846 7857
rect 3790 7783 3846 7792
rect 3712 7670 3832 7698
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3620 5234 3648 7346
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3436 4826 3464 5170
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 3160 3602 3188 3946
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3436 3194 3464 4558
rect 3620 4214 3648 5170
rect 3608 4208 3660 4214
rect 3608 4150 3660 4156
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3528 3534 3556 4082
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3712 3194 3740 7278
rect 3804 4826 3832 7670
rect 3896 6186 3924 11086
rect 3988 10674 4016 11852
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 3988 8090 4016 9658
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4080 6730 4108 11698
rect 4213 10908 4521 10928
rect 4213 10906 4219 10908
rect 4275 10906 4299 10908
rect 4355 10906 4379 10908
rect 4435 10906 4459 10908
rect 4515 10906 4521 10908
rect 4275 10854 4277 10906
rect 4457 10854 4459 10906
rect 4213 10852 4219 10854
rect 4275 10852 4299 10854
rect 4355 10852 4379 10854
rect 4435 10852 4459 10854
rect 4515 10852 4521 10854
rect 4213 10832 4521 10852
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4213 9820 4521 9840
rect 4213 9818 4219 9820
rect 4275 9818 4299 9820
rect 4355 9818 4379 9820
rect 4435 9818 4459 9820
rect 4515 9818 4521 9820
rect 4275 9766 4277 9818
rect 4457 9766 4459 9818
rect 4213 9764 4219 9766
rect 4275 9764 4299 9766
rect 4355 9764 4379 9766
rect 4435 9764 4459 9766
rect 4515 9764 4521 9766
rect 4213 9744 4521 9764
rect 4632 9586 4660 9998
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4213 8732 4521 8752
rect 4213 8730 4219 8732
rect 4275 8730 4299 8732
rect 4355 8730 4379 8732
rect 4435 8730 4459 8732
rect 4515 8730 4521 8732
rect 4275 8678 4277 8730
rect 4457 8678 4459 8730
rect 4213 8676 4219 8678
rect 4275 8676 4299 8678
rect 4355 8676 4379 8678
rect 4435 8676 4459 8678
rect 4515 8676 4521 8678
rect 4213 8656 4521 8676
rect 4213 7644 4521 7664
rect 4213 7642 4219 7644
rect 4275 7642 4299 7644
rect 4355 7642 4379 7644
rect 4435 7642 4459 7644
rect 4515 7642 4521 7644
rect 4275 7590 4277 7642
rect 4457 7590 4459 7642
rect 4213 7588 4219 7590
rect 4275 7588 4299 7590
rect 4355 7588 4379 7590
rect 4435 7588 4459 7590
rect 4515 7588 4521 7590
rect 4213 7568 4521 7588
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4213 6556 4521 6576
rect 4213 6554 4219 6556
rect 4275 6554 4299 6556
rect 4355 6554 4379 6556
rect 4435 6554 4459 6556
rect 4515 6554 4521 6556
rect 4275 6502 4277 6554
rect 4457 6502 4459 6554
rect 4213 6500 4219 6502
rect 4275 6500 4299 6502
rect 4355 6500 4379 6502
rect 4435 6500 4459 6502
rect 4515 6500 4521 6502
rect 4213 6480 4521 6500
rect 3884 6180 3936 6186
rect 3884 6122 3936 6128
rect 4213 5468 4521 5488
rect 4213 5466 4219 5468
rect 4275 5466 4299 5468
rect 4355 5466 4379 5468
rect 4435 5466 4459 5468
rect 4515 5466 4521 5468
rect 4275 5414 4277 5466
rect 4457 5414 4459 5466
rect 4213 5412 4219 5414
rect 4275 5412 4299 5414
rect 4355 5412 4379 5414
rect 4435 5412 4459 5414
rect 4515 5412 4521 5414
rect 4213 5392 4521 5412
rect 4724 5166 4752 29514
rect 5092 29238 5120 42463
rect 5080 29232 5132 29238
rect 5080 29174 5132 29180
rect 5184 27470 5212 45455
rect 5276 32026 5304 56238
rect 5368 46374 5396 57190
rect 5448 54596 5500 54602
rect 5448 54538 5500 54544
rect 5356 46368 5408 46374
rect 5356 46310 5408 46316
rect 5356 46096 5408 46102
rect 5356 46038 5408 46044
rect 5368 45778 5396 46038
rect 5460 45898 5488 54538
rect 5552 48346 5580 76842
rect 5845 76732 6153 76752
rect 5845 76730 5851 76732
rect 5907 76730 5931 76732
rect 5987 76730 6011 76732
rect 6067 76730 6091 76732
rect 6147 76730 6153 76732
rect 5907 76678 5909 76730
rect 6089 76678 6091 76730
rect 5845 76676 5851 76678
rect 5907 76676 5931 76678
rect 5987 76676 6011 76678
rect 6067 76676 6091 76678
rect 6147 76676 6153 76678
rect 5845 76656 6153 76676
rect 9109 76732 9417 76752
rect 9109 76730 9115 76732
rect 9171 76730 9195 76732
rect 9251 76730 9275 76732
rect 9331 76730 9355 76732
rect 9411 76730 9417 76732
rect 9171 76678 9173 76730
rect 9353 76678 9355 76730
rect 9109 76676 9115 76678
rect 9171 76676 9195 76678
rect 9251 76676 9275 76678
rect 9331 76676 9355 76678
rect 9411 76676 9417 76678
rect 9109 76656 9417 76676
rect 10140 76424 10192 76430
rect 10138 76392 10140 76401
rect 10192 76392 10194 76401
rect 10138 76327 10194 76336
rect 9956 76288 10008 76294
rect 9956 76230 10008 76236
rect 7477 76188 7785 76208
rect 7477 76186 7483 76188
rect 7539 76186 7563 76188
rect 7619 76186 7643 76188
rect 7699 76186 7723 76188
rect 7779 76186 7785 76188
rect 7539 76134 7541 76186
rect 7721 76134 7723 76186
rect 7477 76132 7483 76134
rect 7539 76132 7563 76134
rect 7619 76132 7643 76134
rect 7699 76132 7723 76134
rect 7779 76132 7785 76134
rect 7477 76112 7785 76132
rect 5845 75644 6153 75664
rect 5845 75642 5851 75644
rect 5907 75642 5931 75644
rect 5987 75642 6011 75644
rect 6067 75642 6091 75644
rect 6147 75642 6153 75644
rect 5907 75590 5909 75642
rect 6089 75590 6091 75642
rect 5845 75588 5851 75590
rect 5907 75588 5931 75590
rect 5987 75588 6011 75590
rect 6067 75588 6091 75590
rect 6147 75588 6153 75590
rect 5845 75568 6153 75588
rect 9109 75644 9417 75664
rect 9109 75642 9115 75644
rect 9171 75642 9195 75644
rect 9251 75642 9275 75644
rect 9331 75642 9355 75644
rect 9411 75642 9417 75644
rect 9171 75590 9173 75642
rect 9353 75590 9355 75642
rect 9109 75588 9115 75590
rect 9171 75588 9195 75590
rect 9251 75588 9275 75590
rect 9331 75588 9355 75590
rect 9411 75588 9417 75590
rect 9109 75568 9417 75588
rect 8300 75472 8352 75478
rect 8300 75414 8352 75420
rect 7477 75100 7785 75120
rect 7477 75098 7483 75100
rect 7539 75098 7563 75100
rect 7619 75098 7643 75100
rect 7699 75098 7723 75100
rect 7779 75098 7785 75100
rect 7539 75046 7541 75098
rect 7721 75046 7723 75098
rect 7477 75044 7483 75046
rect 7539 75044 7563 75046
rect 7619 75044 7643 75046
rect 7699 75044 7723 75046
rect 7779 75044 7785 75046
rect 7477 75024 7785 75044
rect 5632 74656 5684 74662
rect 5632 74598 5684 74604
rect 5540 48340 5592 48346
rect 5540 48282 5592 48288
rect 5448 45892 5500 45898
rect 5448 45834 5500 45840
rect 5368 45750 5488 45778
rect 5356 45620 5408 45626
rect 5356 45562 5408 45568
rect 5264 32020 5316 32026
rect 5264 31962 5316 31968
rect 5368 30326 5396 45562
rect 5460 35018 5488 45750
rect 5644 45370 5672 74598
rect 5845 74556 6153 74576
rect 5845 74554 5851 74556
rect 5907 74554 5931 74556
rect 5987 74554 6011 74556
rect 6067 74554 6091 74556
rect 6147 74554 6153 74556
rect 5907 74502 5909 74554
rect 6089 74502 6091 74554
rect 5845 74500 5851 74502
rect 5907 74500 5931 74502
rect 5987 74500 6011 74502
rect 6067 74500 6091 74502
rect 6147 74500 6153 74502
rect 5845 74480 6153 74500
rect 7477 74012 7785 74032
rect 7477 74010 7483 74012
rect 7539 74010 7563 74012
rect 7619 74010 7643 74012
rect 7699 74010 7723 74012
rect 7779 74010 7785 74012
rect 7539 73958 7541 74010
rect 7721 73958 7723 74010
rect 7477 73956 7483 73958
rect 7539 73956 7563 73958
rect 7619 73956 7643 73958
rect 7699 73956 7723 73958
rect 7779 73956 7785 73958
rect 7477 73936 7785 73956
rect 5845 73468 6153 73488
rect 5845 73466 5851 73468
rect 5907 73466 5931 73468
rect 5987 73466 6011 73468
rect 6067 73466 6091 73468
rect 6147 73466 6153 73468
rect 5907 73414 5909 73466
rect 6089 73414 6091 73466
rect 5845 73412 5851 73414
rect 5907 73412 5931 73414
rect 5987 73412 6011 73414
rect 6067 73412 6091 73414
rect 6147 73412 6153 73414
rect 5845 73392 6153 73412
rect 7477 72924 7785 72944
rect 7477 72922 7483 72924
rect 7539 72922 7563 72924
rect 7619 72922 7643 72924
rect 7699 72922 7723 72924
rect 7779 72922 7785 72924
rect 7539 72870 7541 72922
rect 7721 72870 7723 72922
rect 7477 72868 7483 72870
rect 7539 72868 7563 72870
rect 7619 72868 7643 72870
rect 7699 72868 7723 72870
rect 7779 72868 7785 72870
rect 7477 72848 7785 72868
rect 5845 72380 6153 72400
rect 5845 72378 5851 72380
rect 5907 72378 5931 72380
rect 5987 72378 6011 72380
rect 6067 72378 6091 72380
rect 6147 72378 6153 72380
rect 5907 72326 5909 72378
rect 6089 72326 6091 72378
rect 5845 72324 5851 72326
rect 5907 72324 5931 72326
rect 5987 72324 6011 72326
rect 6067 72324 6091 72326
rect 6147 72324 6153 72326
rect 5845 72304 6153 72324
rect 7477 71836 7785 71856
rect 7477 71834 7483 71836
rect 7539 71834 7563 71836
rect 7619 71834 7643 71836
rect 7699 71834 7723 71836
rect 7779 71834 7785 71836
rect 7539 71782 7541 71834
rect 7721 71782 7723 71834
rect 7477 71780 7483 71782
rect 7539 71780 7563 71782
rect 7619 71780 7643 71782
rect 7699 71780 7723 71782
rect 7779 71780 7785 71782
rect 7477 71760 7785 71780
rect 5845 71292 6153 71312
rect 5845 71290 5851 71292
rect 5907 71290 5931 71292
rect 5987 71290 6011 71292
rect 6067 71290 6091 71292
rect 6147 71290 6153 71292
rect 5907 71238 5909 71290
rect 6089 71238 6091 71290
rect 5845 71236 5851 71238
rect 5907 71236 5931 71238
rect 5987 71236 6011 71238
rect 6067 71236 6091 71238
rect 6147 71236 6153 71238
rect 5845 71216 6153 71236
rect 7477 70748 7785 70768
rect 7477 70746 7483 70748
rect 7539 70746 7563 70748
rect 7619 70746 7643 70748
rect 7699 70746 7723 70748
rect 7779 70746 7785 70748
rect 7539 70694 7541 70746
rect 7721 70694 7723 70746
rect 7477 70692 7483 70694
rect 7539 70692 7563 70694
rect 7619 70692 7643 70694
rect 7699 70692 7723 70694
rect 7779 70692 7785 70694
rect 7477 70672 7785 70692
rect 5724 70440 5776 70446
rect 5724 70382 5776 70388
rect 5552 45342 5672 45370
rect 5552 44266 5580 45342
rect 5632 45280 5684 45286
rect 5632 45222 5684 45228
rect 5540 44260 5592 44266
rect 5540 44202 5592 44208
rect 5540 43988 5592 43994
rect 5540 43930 5592 43936
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 5356 30320 5408 30326
rect 5356 30262 5408 30268
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 4804 21956 4856 21962
rect 4804 21898 4856 21904
rect 4816 21622 4844 21898
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 5552 5370 5580 43930
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4826 4200 4966
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4724 4758 4752 5102
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2424 2582 2452 2994
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 1400 2440 1452 2446
rect 1400 2382 1452 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2792 649 2820 2382
rect 2884 1465 2912 2382
rect 3620 2281 3648 2994
rect 3804 2650 3832 4490
rect 3988 4457 4016 4558
rect 3974 4448 4030 4457
rect 3974 4383 4030 4392
rect 4213 4380 4521 4400
rect 4213 4378 4219 4380
rect 4275 4378 4299 4380
rect 4355 4378 4379 4380
rect 4435 4378 4459 4380
rect 4515 4378 4521 4380
rect 4275 4326 4277 4378
rect 4457 4326 4459 4378
rect 4213 4324 4219 4326
rect 4275 4324 4299 4326
rect 4355 4324 4379 4326
rect 4435 4324 4459 4326
rect 4515 4324 4521 4326
rect 4213 4304 4521 4324
rect 4620 4072 4672 4078
rect 3974 4040 4030 4049
rect 4620 4014 4672 4020
rect 3974 3975 4030 3984
rect 3988 3534 4016 3975
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 4213 3292 4521 3312
rect 4213 3290 4219 3292
rect 4275 3290 4299 3292
rect 4355 3290 4379 3292
rect 4435 3290 4459 3292
rect 4515 3290 4521 3292
rect 4275 3238 4277 3290
rect 4457 3238 4459 3290
rect 4213 3236 4219 3238
rect 4275 3236 4299 3238
rect 4355 3236 4379 3238
rect 4435 3236 4459 3238
rect 4515 3236 4521 3238
rect 4213 3216 4521 3236
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4066 2544 4122 2553
rect 4172 2530 4200 2994
rect 4632 2650 4660 4014
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5092 2650 5120 2926
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4122 2502 4200 2530
rect 4066 2479 4122 2488
rect 5552 2446 5580 3946
rect 5644 2854 5672 45222
rect 5736 41478 5764 70382
rect 5845 70204 6153 70224
rect 5845 70202 5851 70204
rect 5907 70202 5931 70204
rect 5987 70202 6011 70204
rect 6067 70202 6091 70204
rect 6147 70202 6153 70204
rect 5907 70150 5909 70202
rect 6089 70150 6091 70202
rect 5845 70148 5851 70150
rect 5907 70148 5931 70150
rect 5987 70148 6011 70150
rect 6067 70148 6091 70150
rect 6147 70148 6153 70150
rect 5845 70128 6153 70148
rect 7477 69660 7785 69680
rect 7477 69658 7483 69660
rect 7539 69658 7563 69660
rect 7619 69658 7643 69660
rect 7699 69658 7723 69660
rect 7779 69658 7785 69660
rect 7539 69606 7541 69658
rect 7721 69606 7723 69658
rect 7477 69604 7483 69606
rect 7539 69604 7563 69606
rect 7619 69604 7643 69606
rect 7699 69604 7723 69606
rect 7779 69604 7785 69606
rect 7477 69584 7785 69604
rect 5845 69116 6153 69136
rect 5845 69114 5851 69116
rect 5907 69114 5931 69116
rect 5987 69114 6011 69116
rect 6067 69114 6091 69116
rect 6147 69114 6153 69116
rect 5907 69062 5909 69114
rect 6089 69062 6091 69114
rect 5845 69060 5851 69062
rect 5907 69060 5931 69062
rect 5987 69060 6011 69062
rect 6067 69060 6091 69062
rect 6147 69060 6153 69062
rect 5845 69040 6153 69060
rect 7012 68672 7064 68678
rect 7012 68614 7064 68620
rect 5845 68028 6153 68048
rect 5845 68026 5851 68028
rect 5907 68026 5931 68028
rect 5987 68026 6011 68028
rect 6067 68026 6091 68028
rect 6147 68026 6153 68028
rect 5907 67974 5909 68026
rect 6089 67974 6091 68026
rect 5845 67972 5851 67974
rect 5907 67972 5931 67974
rect 5987 67972 6011 67974
rect 6067 67972 6091 67974
rect 6147 67972 6153 67974
rect 5845 67952 6153 67972
rect 5845 66940 6153 66960
rect 5845 66938 5851 66940
rect 5907 66938 5931 66940
rect 5987 66938 6011 66940
rect 6067 66938 6091 66940
rect 6147 66938 6153 66940
rect 5907 66886 5909 66938
rect 6089 66886 6091 66938
rect 5845 66884 5851 66886
rect 5907 66884 5931 66886
rect 5987 66884 6011 66886
rect 6067 66884 6091 66886
rect 6147 66884 6153 66886
rect 5845 66864 6153 66884
rect 5845 65852 6153 65872
rect 5845 65850 5851 65852
rect 5907 65850 5931 65852
rect 5987 65850 6011 65852
rect 6067 65850 6091 65852
rect 6147 65850 6153 65852
rect 5907 65798 5909 65850
rect 6089 65798 6091 65850
rect 5845 65796 5851 65798
rect 5907 65796 5931 65798
rect 5987 65796 6011 65798
rect 6067 65796 6091 65798
rect 6147 65796 6153 65798
rect 5845 65776 6153 65796
rect 5908 65680 5960 65686
rect 5906 65648 5908 65657
rect 5960 65648 5962 65657
rect 5906 65583 5962 65592
rect 6828 65204 6880 65210
rect 6828 65146 6880 65152
rect 6368 64864 6420 64870
rect 6368 64806 6420 64812
rect 5845 64764 6153 64784
rect 5845 64762 5851 64764
rect 5907 64762 5931 64764
rect 5987 64762 6011 64764
rect 6067 64762 6091 64764
rect 6147 64762 6153 64764
rect 5907 64710 5909 64762
rect 6089 64710 6091 64762
rect 5845 64708 5851 64710
rect 5907 64708 5931 64710
rect 5987 64708 6011 64710
rect 6067 64708 6091 64710
rect 6147 64708 6153 64710
rect 5845 64688 6153 64708
rect 6380 64394 6408 64806
rect 6368 64388 6420 64394
rect 6368 64330 6420 64336
rect 5845 63676 6153 63696
rect 5845 63674 5851 63676
rect 5907 63674 5931 63676
rect 5987 63674 6011 63676
rect 6067 63674 6091 63676
rect 6147 63674 6153 63676
rect 5907 63622 5909 63674
rect 6089 63622 6091 63674
rect 5845 63620 5851 63622
rect 5907 63620 5931 63622
rect 5987 63620 6011 63622
rect 6067 63620 6091 63622
rect 6147 63620 6153 63622
rect 5845 63600 6153 63620
rect 5845 62588 6153 62608
rect 5845 62586 5851 62588
rect 5907 62586 5931 62588
rect 5987 62586 6011 62588
rect 6067 62586 6091 62588
rect 6147 62586 6153 62588
rect 5907 62534 5909 62586
rect 6089 62534 6091 62586
rect 5845 62532 5851 62534
rect 5907 62532 5931 62534
rect 5987 62532 6011 62534
rect 6067 62532 6091 62534
rect 6147 62532 6153 62534
rect 5845 62512 6153 62532
rect 5845 61500 6153 61520
rect 5845 61498 5851 61500
rect 5907 61498 5931 61500
rect 5987 61498 6011 61500
rect 6067 61498 6091 61500
rect 6147 61498 6153 61500
rect 5907 61446 5909 61498
rect 6089 61446 6091 61498
rect 5845 61444 5851 61446
rect 5907 61444 5931 61446
rect 5987 61444 6011 61446
rect 6067 61444 6091 61446
rect 6147 61444 6153 61446
rect 5845 61424 6153 61444
rect 6368 60512 6420 60518
rect 6368 60454 6420 60460
rect 5845 60412 6153 60432
rect 5845 60410 5851 60412
rect 5907 60410 5931 60412
rect 5987 60410 6011 60412
rect 6067 60410 6091 60412
rect 6147 60410 6153 60412
rect 5907 60358 5909 60410
rect 6089 60358 6091 60410
rect 5845 60356 5851 60358
rect 5907 60356 5931 60358
rect 5987 60356 6011 60358
rect 6067 60356 6091 60358
rect 6147 60356 6153 60358
rect 5845 60336 6153 60356
rect 5845 59324 6153 59344
rect 5845 59322 5851 59324
rect 5907 59322 5931 59324
rect 5987 59322 6011 59324
rect 6067 59322 6091 59324
rect 6147 59322 6153 59324
rect 5907 59270 5909 59322
rect 6089 59270 6091 59322
rect 5845 59268 5851 59270
rect 5907 59268 5931 59270
rect 5987 59268 6011 59270
rect 6067 59268 6091 59270
rect 6147 59268 6153 59270
rect 5845 59248 6153 59268
rect 5845 58236 6153 58256
rect 5845 58234 5851 58236
rect 5907 58234 5931 58236
rect 5987 58234 6011 58236
rect 6067 58234 6091 58236
rect 6147 58234 6153 58236
rect 5907 58182 5909 58234
rect 6089 58182 6091 58234
rect 5845 58180 5851 58182
rect 5907 58180 5931 58182
rect 5987 58180 6011 58182
rect 6067 58180 6091 58182
rect 6147 58180 6153 58182
rect 5845 58160 6153 58180
rect 5845 57148 6153 57168
rect 5845 57146 5851 57148
rect 5907 57146 5931 57148
rect 5987 57146 6011 57148
rect 6067 57146 6091 57148
rect 6147 57146 6153 57148
rect 5907 57094 5909 57146
rect 6089 57094 6091 57146
rect 5845 57092 5851 57094
rect 5907 57092 5931 57094
rect 5987 57092 6011 57094
rect 6067 57092 6091 57094
rect 6147 57092 6153 57094
rect 5845 57072 6153 57092
rect 5845 56060 6153 56080
rect 5845 56058 5851 56060
rect 5907 56058 5931 56060
rect 5987 56058 6011 56060
rect 6067 56058 6091 56060
rect 6147 56058 6153 56060
rect 5907 56006 5909 56058
rect 6089 56006 6091 56058
rect 5845 56004 5851 56006
rect 5907 56004 5931 56006
rect 5987 56004 6011 56006
rect 6067 56004 6091 56006
rect 6147 56004 6153 56006
rect 5845 55984 6153 56004
rect 5845 54972 6153 54992
rect 5845 54970 5851 54972
rect 5907 54970 5931 54972
rect 5987 54970 6011 54972
rect 6067 54970 6091 54972
rect 6147 54970 6153 54972
rect 5907 54918 5909 54970
rect 6089 54918 6091 54970
rect 5845 54916 5851 54918
rect 5907 54916 5931 54918
rect 5987 54916 6011 54918
rect 6067 54916 6091 54918
rect 6147 54916 6153 54918
rect 5845 54896 6153 54916
rect 5845 53884 6153 53904
rect 5845 53882 5851 53884
rect 5907 53882 5931 53884
rect 5987 53882 6011 53884
rect 6067 53882 6091 53884
rect 6147 53882 6153 53884
rect 5907 53830 5909 53882
rect 6089 53830 6091 53882
rect 5845 53828 5851 53830
rect 5907 53828 5931 53830
rect 5987 53828 6011 53830
rect 6067 53828 6091 53830
rect 6147 53828 6153 53830
rect 5845 53808 6153 53828
rect 5845 52796 6153 52816
rect 5845 52794 5851 52796
rect 5907 52794 5931 52796
rect 5987 52794 6011 52796
rect 6067 52794 6091 52796
rect 6147 52794 6153 52796
rect 5907 52742 5909 52794
rect 6089 52742 6091 52794
rect 5845 52740 5851 52742
rect 5907 52740 5931 52742
rect 5987 52740 6011 52742
rect 6067 52740 6091 52742
rect 6147 52740 6153 52742
rect 5845 52720 6153 52740
rect 6276 52624 6328 52630
rect 6276 52566 6328 52572
rect 5845 51708 6153 51728
rect 5845 51706 5851 51708
rect 5907 51706 5931 51708
rect 5987 51706 6011 51708
rect 6067 51706 6091 51708
rect 6147 51706 6153 51708
rect 5907 51654 5909 51706
rect 6089 51654 6091 51706
rect 5845 51652 5851 51654
rect 5907 51652 5931 51654
rect 5987 51652 6011 51654
rect 6067 51652 6091 51654
rect 6147 51652 6153 51654
rect 5845 51632 6153 51652
rect 5845 50620 6153 50640
rect 5845 50618 5851 50620
rect 5907 50618 5931 50620
rect 5987 50618 6011 50620
rect 6067 50618 6091 50620
rect 6147 50618 6153 50620
rect 5907 50566 5909 50618
rect 6089 50566 6091 50618
rect 5845 50564 5851 50566
rect 5907 50564 5931 50566
rect 5987 50564 6011 50566
rect 6067 50564 6091 50566
rect 6147 50564 6153 50566
rect 5845 50544 6153 50564
rect 6184 49836 6236 49842
rect 6184 49778 6236 49784
rect 5845 49532 6153 49552
rect 5845 49530 5851 49532
rect 5907 49530 5931 49532
rect 5987 49530 6011 49532
rect 6067 49530 6091 49532
rect 6147 49530 6153 49532
rect 5907 49478 5909 49530
rect 6089 49478 6091 49530
rect 5845 49476 5851 49478
rect 5907 49476 5931 49478
rect 5987 49476 6011 49478
rect 6067 49476 6091 49478
rect 6147 49476 6153 49478
rect 5845 49456 6153 49476
rect 5845 48444 6153 48464
rect 5845 48442 5851 48444
rect 5907 48442 5931 48444
rect 5987 48442 6011 48444
rect 6067 48442 6091 48444
rect 6147 48442 6153 48444
rect 5907 48390 5909 48442
rect 6089 48390 6091 48442
rect 5845 48388 5851 48390
rect 5907 48388 5931 48390
rect 5987 48388 6011 48390
rect 6067 48388 6091 48390
rect 6147 48388 6153 48390
rect 5845 48368 6153 48388
rect 6196 48328 6224 49778
rect 5920 48300 6224 48328
rect 5920 47569 5948 48300
rect 6184 48068 6236 48074
rect 6184 48010 6236 48016
rect 5906 47560 5962 47569
rect 5906 47495 5962 47504
rect 5845 47356 6153 47376
rect 5845 47354 5851 47356
rect 5907 47354 5931 47356
rect 5987 47354 6011 47356
rect 6067 47354 6091 47356
rect 6147 47354 6153 47356
rect 5907 47302 5909 47354
rect 6089 47302 6091 47354
rect 5845 47300 5851 47302
rect 5907 47300 5931 47302
rect 5987 47300 6011 47302
rect 6067 47300 6091 47302
rect 6147 47300 6153 47302
rect 5845 47280 6153 47300
rect 5845 46268 6153 46288
rect 5845 46266 5851 46268
rect 5907 46266 5931 46268
rect 5987 46266 6011 46268
rect 6067 46266 6091 46268
rect 6147 46266 6153 46268
rect 5907 46214 5909 46266
rect 6089 46214 6091 46266
rect 5845 46212 5851 46214
rect 5907 46212 5931 46214
rect 5987 46212 6011 46214
rect 6067 46212 6091 46214
rect 6147 46212 6153 46214
rect 5845 46192 6153 46212
rect 5845 45180 6153 45200
rect 5845 45178 5851 45180
rect 5907 45178 5931 45180
rect 5987 45178 6011 45180
rect 6067 45178 6091 45180
rect 6147 45178 6153 45180
rect 5907 45126 5909 45178
rect 6089 45126 6091 45178
rect 5845 45124 5851 45126
rect 5907 45124 5931 45126
rect 5987 45124 6011 45126
rect 6067 45124 6091 45126
rect 6147 45124 6153 45126
rect 5845 45104 6153 45124
rect 5845 44092 6153 44112
rect 5845 44090 5851 44092
rect 5907 44090 5931 44092
rect 5987 44090 6011 44092
rect 6067 44090 6091 44092
rect 6147 44090 6153 44092
rect 5907 44038 5909 44090
rect 6089 44038 6091 44090
rect 5845 44036 5851 44038
rect 5907 44036 5931 44038
rect 5987 44036 6011 44038
rect 6067 44036 6091 44038
rect 6147 44036 6153 44038
rect 5845 44016 6153 44036
rect 6196 43994 6224 48010
rect 6184 43988 6236 43994
rect 6184 43930 6236 43936
rect 6184 43852 6236 43858
rect 6184 43794 6236 43800
rect 5845 43004 6153 43024
rect 5845 43002 5851 43004
rect 5907 43002 5931 43004
rect 5987 43002 6011 43004
rect 6067 43002 6091 43004
rect 6147 43002 6153 43004
rect 5907 42950 5909 43002
rect 6089 42950 6091 43002
rect 5845 42948 5851 42950
rect 5907 42948 5931 42950
rect 5987 42948 6011 42950
rect 6067 42948 6091 42950
rect 6147 42948 6153 42950
rect 5845 42928 6153 42948
rect 5845 41916 6153 41936
rect 5845 41914 5851 41916
rect 5907 41914 5931 41916
rect 5987 41914 6011 41916
rect 6067 41914 6091 41916
rect 6147 41914 6153 41916
rect 5907 41862 5909 41914
rect 6089 41862 6091 41914
rect 5845 41860 5851 41862
rect 5907 41860 5931 41862
rect 5987 41860 6011 41862
rect 6067 41860 6091 41862
rect 6147 41860 6153 41862
rect 5845 41840 6153 41860
rect 5724 41472 5776 41478
rect 5724 41414 5776 41420
rect 5845 40828 6153 40848
rect 5845 40826 5851 40828
rect 5907 40826 5931 40828
rect 5987 40826 6011 40828
rect 6067 40826 6091 40828
rect 6147 40826 6153 40828
rect 5907 40774 5909 40826
rect 6089 40774 6091 40826
rect 5845 40772 5851 40774
rect 5907 40772 5931 40774
rect 5987 40772 6011 40774
rect 6067 40772 6091 40774
rect 6147 40772 6153 40774
rect 5845 40752 6153 40772
rect 5845 39740 6153 39760
rect 5845 39738 5851 39740
rect 5907 39738 5931 39740
rect 5987 39738 6011 39740
rect 6067 39738 6091 39740
rect 6147 39738 6153 39740
rect 5907 39686 5909 39738
rect 6089 39686 6091 39738
rect 5845 39684 5851 39686
rect 5907 39684 5931 39686
rect 5987 39684 6011 39686
rect 6067 39684 6091 39686
rect 6147 39684 6153 39686
rect 5845 39664 6153 39684
rect 5845 38652 6153 38672
rect 5845 38650 5851 38652
rect 5907 38650 5931 38652
rect 5987 38650 6011 38652
rect 6067 38650 6091 38652
rect 6147 38650 6153 38652
rect 5907 38598 5909 38650
rect 6089 38598 6091 38650
rect 5845 38596 5851 38598
rect 5907 38596 5931 38598
rect 5987 38596 6011 38598
rect 6067 38596 6091 38598
rect 6147 38596 6153 38598
rect 5845 38576 6153 38596
rect 5845 37564 6153 37584
rect 5845 37562 5851 37564
rect 5907 37562 5931 37564
rect 5987 37562 6011 37564
rect 6067 37562 6091 37564
rect 6147 37562 6153 37564
rect 5907 37510 5909 37562
rect 6089 37510 6091 37562
rect 5845 37508 5851 37510
rect 5907 37508 5931 37510
rect 5987 37508 6011 37510
rect 6067 37508 6091 37510
rect 6147 37508 6153 37510
rect 5845 37488 6153 37508
rect 5845 36476 6153 36496
rect 5845 36474 5851 36476
rect 5907 36474 5931 36476
rect 5987 36474 6011 36476
rect 6067 36474 6091 36476
rect 6147 36474 6153 36476
rect 5907 36422 5909 36474
rect 6089 36422 6091 36474
rect 5845 36420 5851 36422
rect 5907 36420 5931 36422
rect 5987 36420 6011 36422
rect 6067 36420 6091 36422
rect 6147 36420 6153 36422
rect 5845 36400 6153 36420
rect 5845 35388 6153 35408
rect 5845 35386 5851 35388
rect 5907 35386 5931 35388
rect 5987 35386 6011 35388
rect 6067 35386 6091 35388
rect 6147 35386 6153 35388
rect 5907 35334 5909 35386
rect 6089 35334 6091 35386
rect 5845 35332 5851 35334
rect 5907 35332 5931 35334
rect 5987 35332 6011 35334
rect 6067 35332 6091 35334
rect 6147 35332 6153 35334
rect 5845 35312 6153 35332
rect 5845 34300 6153 34320
rect 5845 34298 5851 34300
rect 5907 34298 5931 34300
rect 5987 34298 6011 34300
rect 6067 34298 6091 34300
rect 6147 34298 6153 34300
rect 5907 34246 5909 34298
rect 6089 34246 6091 34298
rect 5845 34244 5851 34246
rect 5907 34244 5931 34246
rect 5987 34244 6011 34246
rect 6067 34244 6091 34246
rect 6147 34244 6153 34246
rect 5845 34224 6153 34244
rect 5845 33212 6153 33232
rect 5845 33210 5851 33212
rect 5907 33210 5931 33212
rect 5987 33210 6011 33212
rect 6067 33210 6091 33212
rect 6147 33210 6153 33212
rect 5907 33158 5909 33210
rect 6089 33158 6091 33210
rect 5845 33156 5851 33158
rect 5907 33156 5931 33158
rect 5987 33156 6011 33158
rect 6067 33156 6091 33158
rect 6147 33156 6153 33158
rect 5845 33136 6153 33156
rect 5845 32124 6153 32144
rect 5845 32122 5851 32124
rect 5907 32122 5931 32124
rect 5987 32122 6011 32124
rect 6067 32122 6091 32124
rect 6147 32122 6153 32124
rect 5907 32070 5909 32122
rect 6089 32070 6091 32122
rect 5845 32068 5851 32070
rect 5907 32068 5931 32070
rect 5987 32068 6011 32070
rect 6067 32068 6091 32070
rect 6147 32068 6153 32070
rect 5845 32048 6153 32068
rect 5845 31036 6153 31056
rect 5845 31034 5851 31036
rect 5907 31034 5931 31036
rect 5987 31034 6011 31036
rect 6067 31034 6091 31036
rect 6147 31034 6153 31036
rect 5907 30982 5909 31034
rect 6089 30982 6091 31034
rect 5845 30980 5851 30982
rect 5907 30980 5931 30982
rect 5987 30980 6011 30982
rect 6067 30980 6091 30982
rect 6147 30980 6153 30982
rect 5845 30960 6153 30980
rect 5845 29948 6153 29968
rect 5845 29946 5851 29948
rect 5907 29946 5931 29948
rect 5987 29946 6011 29948
rect 6067 29946 6091 29948
rect 6147 29946 6153 29948
rect 5907 29894 5909 29946
rect 6089 29894 6091 29946
rect 5845 29892 5851 29894
rect 5907 29892 5931 29894
rect 5987 29892 6011 29894
rect 6067 29892 6091 29894
rect 6147 29892 6153 29894
rect 5845 29872 6153 29892
rect 5845 28860 6153 28880
rect 5845 28858 5851 28860
rect 5907 28858 5931 28860
rect 5987 28858 6011 28860
rect 6067 28858 6091 28860
rect 6147 28858 6153 28860
rect 5907 28806 5909 28858
rect 6089 28806 6091 28858
rect 5845 28804 5851 28806
rect 5907 28804 5931 28806
rect 5987 28804 6011 28806
rect 6067 28804 6091 28806
rect 6147 28804 6153 28806
rect 5845 28784 6153 28804
rect 5845 27772 6153 27792
rect 5845 27770 5851 27772
rect 5907 27770 5931 27772
rect 5987 27770 6011 27772
rect 6067 27770 6091 27772
rect 6147 27770 6153 27772
rect 5907 27718 5909 27770
rect 6089 27718 6091 27770
rect 5845 27716 5851 27718
rect 5907 27716 5931 27718
rect 5987 27716 6011 27718
rect 6067 27716 6091 27718
rect 6147 27716 6153 27718
rect 5845 27696 6153 27716
rect 5845 26684 6153 26704
rect 5845 26682 5851 26684
rect 5907 26682 5931 26684
rect 5987 26682 6011 26684
rect 6067 26682 6091 26684
rect 6147 26682 6153 26684
rect 5907 26630 5909 26682
rect 6089 26630 6091 26682
rect 5845 26628 5851 26630
rect 5907 26628 5931 26630
rect 5987 26628 6011 26630
rect 6067 26628 6091 26630
rect 6147 26628 6153 26630
rect 5845 26608 6153 26628
rect 5845 25596 6153 25616
rect 5845 25594 5851 25596
rect 5907 25594 5931 25596
rect 5987 25594 6011 25596
rect 6067 25594 6091 25596
rect 6147 25594 6153 25596
rect 5907 25542 5909 25594
rect 6089 25542 6091 25594
rect 5845 25540 5851 25542
rect 5907 25540 5931 25542
rect 5987 25540 6011 25542
rect 6067 25540 6091 25542
rect 6147 25540 6153 25542
rect 5845 25520 6153 25540
rect 5845 24508 6153 24528
rect 5845 24506 5851 24508
rect 5907 24506 5931 24508
rect 5987 24506 6011 24508
rect 6067 24506 6091 24508
rect 6147 24506 6153 24508
rect 5907 24454 5909 24506
rect 6089 24454 6091 24506
rect 5845 24452 5851 24454
rect 5907 24452 5931 24454
rect 5987 24452 6011 24454
rect 6067 24452 6091 24454
rect 6147 24452 6153 24454
rect 5845 24432 6153 24452
rect 5845 23420 6153 23440
rect 5845 23418 5851 23420
rect 5907 23418 5931 23420
rect 5987 23418 6011 23420
rect 6067 23418 6091 23420
rect 6147 23418 6153 23420
rect 5907 23366 5909 23418
rect 6089 23366 6091 23418
rect 5845 23364 5851 23366
rect 5907 23364 5931 23366
rect 5987 23364 6011 23366
rect 6067 23364 6091 23366
rect 6147 23364 6153 23366
rect 5845 23344 6153 23364
rect 5845 22332 6153 22352
rect 5845 22330 5851 22332
rect 5907 22330 5931 22332
rect 5987 22330 6011 22332
rect 6067 22330 6091 22332
rect 6147 22330 6153 22332
rect 5907 22278 5909 22330
rect 6089 22278 6091 22330
rect 5845 22276 5851 22278
rect 5907 22276 5931 22278
rect 5987 22276 6011 22278
rect 6067 22276 6091 22278
rect 6147 22276 6153 22278
rect 5845 22256 6153 22276
rect 5845 21244 6153 21264
rect 5845 21242 5851 21244
rect 5907 21242 5931 21244
rect 5987 21242 6011 21244
rect 6067 21242 6091 21244
rect 6147 21242 6153 21244
rect 5907 21190 5909 21242
rect 6089 21190 6091 21242
rect 5845 21188 5851 21190
rect 5907 21188 5931 21190
rect 5987 21188 6011 21190
rect 6067 21188 6091 21190
rect 6147 21188 6153 21190
rect 5845 21168 6153 21188
rect 5845 20156 6153 20176
rect 5845 20154 5851 20156
rect 5907 20154 5931 20156
rect 5987 20154 6011 20156
rect 6067 20154 6091 20156
rect 6147 20154 6153 20156
rect 5907 20102 5909 20154
rect 6089 20102 6091 20154
rect 5845 20100 5851 20102
rect 5907 20100 5931 20102
rect 5987 20100 6011 20102
rect 6067 20100 6091 20102
rect 6147 20100 6153 20102
rect 5845 20080 6153 20100
rect 5845 19068 6153 19088
rect 5845 19066 5851 19068
rect 5907 19066 5931 19068
rect 5987 19066 6011 19068
rect 6067 19066 6091 19068
rect 6147 19066 6153 19068
rect 5907 19014 5909 19066
rect 6089 19014 6091 19066
rect 5845 19012 5851 19014
rect 5907 19012 5931 19014
rect 5987 19012 6011 19014
rect 6067 19012 6091 19014
rect 6147 19012 6153 19014
rect 5845 18992 6153 19012
rect 5845 17980 6153 18000
rect 5845 17978 5851 17980
rect 5907 17978 5931 17980
rect 5987 17978 6011 17980
rect 6067 17978 6091 17980
rect 6147 17978 6153 17980
rect 5907 17926 5909 17978
rect 6089 17926 6091 17978
rect 5845 17924 5851 17926
rect 5907 17924 5931 17926
rect 5987 17924 6011 17926
rect 6067 17924 6091 17926
rect 6147 17924 6153 17926
rect 5845 17904 6153 17924
rect 5845 16892 6153 16912
rect 5845 16890 5851 16892
rect 5907 16890 5931 16892
rect 5987 16890 6011 16892
rect 6067 16890 6091 16892
rect 6147 16890 6153 16892
rect 5907 16838 5909 16890
rect 6089 16838 6091 16890
rect 5845 16836 5851 16838
rect 5907 16836 5931 16838
rect 5987 16836 6011 16838
rect 6067 16836 6091 16838
rect 6147 16836 6153 16838
rect 5845 16816 6153 16836
rect 5845 15804 6153 15824
rect 5845 15802 5851 15804
rect 5907 15802 5931 15804
rect 5987 15802 6011 15804
rect 6067 15802 6091 15804
rect 6147 15802 6153 15804
rect 5907 15750 5909 15802
rect 6089 15750 6091 15802
rect 5845 15748 5851 15750
rect 5907 15748 5931 15750
rect 5987 15748 6011 15750
rect 6067 15748 6091 15750
rect 6147 15748 6153 15750
rect 5845 15728 6153 15748
rect 5845 14716 6153 14736
rect 5845 14714 5851 14716
rect 5907 14714 5931 14716
rect 5987 14714 6011 14716
rect 6067 14714 6091 14716
rect 6147 14714 6153 14716
rect 5907 14662 5909 14714
rect 6089 14662 6091 14714
rect 5845 14660 5851 14662
rect 5907 14660 5931 14662
rect 5987 14660 6011 14662
rect 6067 14660 6091 14662
rect 6147 14660 6153 14662
rect 5845 14640 6153 14660
rect 5845 13628 6153 13648
rect 5845 13626 5851 13628
rect 5907 13626 5931 13628
rect 5987 13626 6011 13628
rect 6067 13626 6091 13628
rect 6147 13626 6153 13628
rect 5907 13574 5909 13626
rect 6089 13574 6091 13626
rect 5845 13572 5851 13574
rect 5907 13572 5931 13574
rect 5987 13572 6011 13574
rect 6067 13572 6091 13574
rect 6147 13572 6153 13574
rect 5845 13552 6153 13572
rect 5845 12540 6153 12560
rect 5845 12538 5851 12540
rect 5907 12538 5931 12540
rect 5987 12538 6011 12540
rect 6067 12538 6091 12540
rect 6147 12538 6153 12540
rect 5907 12486 5909 12538
rect 6089 12486 6091 12538
rect 5845 12484 5851 12486
rect 5907 12484 5931 12486
rect 5987 12484 6011 12486
rect 6067 12484 6091 12486
rect 6147 12484 6153 12486
rect 5845 12464 6153 12484
rect 5845 11452 6153 11472
rect 5845 11450 5851 11452
rect 5907 11450 5931 11452
rect 5987 11450 6011 11452
rect 6067 11450 6091 11452
rect 6147 11450 6153 11452
rect 5907 11398 5909 11450
rect 6089 11398 6091 11450
rect 5845 11396 5851 11398
rect 5907 11396 5931 11398
rect 5987 11396 6011 11398
rect 6067 11396 6091 11398
rect 6147 11396 6153 11398
rect 5845 11376 6153 11396
rect 5845 10364 6153 10384
rect 5845 10362 5851 10364
rect 5907 10362 5931 10364
rect 5987 10362 6011 10364
rect 6067 10362 6091 10364
rect 6147 10362 6153 10364
rect 5907 10310 5909 10362
rect 6089 10310 6091 10362
rect 5845 10308 5851 10310
rect 5907 10308 5931 10310
rect 5987 10308 6011 10310
rect 6067 10308 6091 10310
rect 6147 10308 6153 10310
rect 5845 10288 6153 10308
rect 5845 9276 6153 9296
rect 5845 9274 5851 9276
rect 5907 9274 5931 9276
rect 5987 9274 6011 9276
rect 6067 9274 6091 9276
rect 6147 9274 6153 9276
rect 5907 9222 5909 9274
rect 6089 9222 6091 9274
rect 5845 9220 5851 9222
rect 5907 9220 5931 9222
rect 5987 9220 6011 9222
rect 6067 9220 6091 9222
rect 6147 9220 6153 9222
rect 5845 9200 6153 9220
rect 6196 8838 6224 43794
rect 6288 22710 6316 52566
rect 6380 38758 6408 60454
rect 6644 56908 6696 56914
rect 6644 56850 6696 56856
rect 6552 48748 6604 48754
rect 6552 48690 6604 48696
rect 6460 48680 6512 48686
rect 6460 48622 6512 48628
rect 6368 38752 6420 38758
rect 6368 38694 6420 38700
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 6472 8906 6500 48622
rect 6564 9110 6592 48690
rect 6656 31482 6684 56850
rect 6736 49292 6788 49298
rect 6736 49234 6788 49240
rect 6748 43858 6776 49234
rect 6840 44878 6868 65146
rect 6920 64592 6972 64598
rect 6920 64534 6972 64540
rect 6828 44872 6880 44878
rect 6828 44814 6880 44820
rect 6736 43852 6788 43858
rect 6736 43794 6788 43800
rect 6734 43752 6790 43761
rect 6734 43687 6790 43696
rect 6644 31476 6696 31482
rect 6644 31418 6696 31424
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6748 8566 6776 43687
rect 6932 36854 6960 64534
rect 7024 41682 7052 68614
rect 7477 68572 7785 68592
rect 7477 68570 7483 68572
rect 7539 68570 7563 68572
rect 7619 68570 7643 68572
rect 7699 68570 7723 68572
rect 7779 68570 7785 68572
rect 7539 68518 7541 68570
rect 7721 68518 7723 68570
rect 7477 68516 7483 68518
rect 7539 68516 7563 68518
rect 7619 68516 7643 68518
rect 7699 68516 7723 68518
rect 7779 68516 7785 68518
rect 7477 68496 7785 68516
rect 7477 67484 7785 67504
rect 7477 67482 7483 67484
rect 7539 67482 7563 67484
rect 7619 67482 7643 67484
rect 7699 67482 7723 67484
rect 7779 67482 7785 67484
rect 7539 67430 7541 67482
rect 7721 67430 7723 67482
rect 7477 67428 7483 67430
rect 7539 67428 7563 67430
rect 7619 67428 7643 67430
rect 7699 67428 7723 67430
rect 7779 67428 7785 67430
rect 7477 67408 7785 67428
rect 7477 66396 7785 66416
rect 7477 66394 7483 66396
rect 7539 66394 7563 66396
rect 7619 66394 7643 66396
rect 7699 66394 7723 66396
rect 7779 66394 7785 66396
rect 7539 66342 7541 66394
rect 7721 66342 7723 66394
rect 7477 66340 7483 66342
rect 7539 66340 7563 66342
rect 7619 66340 7643 66342
rect 7699 66340 7723 66342
rect 7779 66340 7785 66342
rect 7477 66320 7785 66340
rect 7194 66192 7250 66201
rect 7194 66127 7250 66136
rect 7208 66026 7236 66127
rect 7104 66020 7156 66026
rect 7104 65962 7156 65968
rect 7196 66020 7248 66026
rect 7196 65962 7248 65968
rect 7116 65754 7144 65962
rect 7104 65748 7156 65754
rect 7104 65690 7156 65696
rect 7477 65308 7785 65328
rect 7477 65306 7483 65308
rect 7539 65306 7563 65308
rect 7619 65306 7643 65308
rect 7699 65306 7723 65308
rect 7779 65306 7785 65308
rect 7539 65254 7541 65306
rect 7721 65254 7723 65306
rect 7477 65252 7483 65254
rect 7539 65252 7563 65254
rect 7619 65252 7643 65254
rect 7699 65252 7723 65254
rect 7779 65252 7785 65254
rect 7477 65232 7785 65252
rect 7477 64220 7785 64240
rect 7477 64218 7483 64220
rect 7539 64218 7563 64220
rect 7619 64218 7643 64220
rect 7699 64218 7723 64220
rect 7779 64218 7785 64220
rect 7539 64166 7541 64218
rect 7721 64166 7723 64218
rect 7477 64164 7483 64166
rect 7539 64164 7563 64166
rect 7619 64164 7643 64166
rect 7699 64164 7723 64166
rect 7779 64164 7785 64166
rect 7477 64144 7785 64164
rect 7477 63132 7785 63152
rect 7477 63130 7483 63132
rect 7539 63130 7563 63132
rect 7619 63130 7643 63132
rect 7699 63130 7723 63132
rect 7779 63130 7785 63132
rect 7539 63078 7541 63130
rect 7721 63078 7723 63130
rect 7477 63076 7483 63078
rect 7539 63076 7563 63078
rect 7619 63076 7643 63078
rect 7699 63076 7723 63078
rect 7779 63076 7785 63078
rect 7477 63056 7785 63076
rect 7477 62044 7785 62064
rect 7477 62042 7483 62044
rect 7539 62042 7563 62044
rect 7619 62042 7643 62044
rect 7699 62042 7723 62044
rect 7779 62042 7785 62044
rect 7539 61990 7541 62042
rect 7721 61990 7723 62042
rect 7477 61988 7483 61990
rect 7539 61988 7563 61990
rect 7619 61988 7643 61990
rect 7699 61988 7723 61990
rect 7779 61988 7785 61990
rect 7477 61968 7785 61988
rect 7477 60956 7785 60976
rect 7477 60954 7483 60956
rect 7539 60954 7563 60956
rect 7619 60954 7643 60956
rect 7699 60954 7723 60956
rect 7779 60954 7785 60956
rect 7539 60902 7541 60954
rect 7721 60902 7723 60954
rect 7477 60900 7483 60902
rect 7539 60900 7563 60902
rect 7619 60900 7643 60902
rect 7699 60900 7723 60902
rect 7779 60900 7785 60902
rect 7477 60880 7785 60900
rect 7477 59868 7785 59888
rect 7477 59866 7483 59868
rect 7539 59866 7563 59868
rect 7619 59866 7643 59868
rect 7699 59866 7723 59868
rect 7779 59866 7785 59868
rect 7539 59814 7541 59866
rect 7721 59814 7723 59866
rect 7477 59812 7483 59814
rect 7539 59812 7563 59814
rect 7619 59812 7643 59814
rect 7699 59812 7723 59814
rect 7779 59812 7785 59814
rect 7477 59792 7785 59812
rect 7477 58780 7785 58800
rect 7477 58778 7483 58780
rect 7539 58778 7563 58780
rect 7619 58778 7643 58780
rect 7699 58778 7723 58780
rect 7779 58778 7785 58780
rect 7539 58726 7541 58778
rect 7721 58726 7723 58778
rect 7477 58724 7483 58726
rect 7539 58724 7563 58726
rect 7619 58724 7643 58726
rect 7699 58724 7723 58726
rect 7779 58724 7785 58726
rect 7477 58704 7785 58724
rect 7477 57692 7785 57712
rect 7477 57690 7483 57692
rect 7539 57690 7563 57692
rect 7619 57690 7643 57692
rect 7699 57690 7723 57692
rect 7779 57690 7785 57692
rect 7539 57638 7541 57690
rect 7721 57638 7723 57690
rect 7477 57636 7483 57638
rect 7539 57636 7563 57638
rect 7619 57636 7643 57638
rect 7699 57636 7723 57638
rect 7779 57636 7785 57638
rect 7477 57616 7785 57636
rect 7477 56604 7785 56624
rect 7477 56602 7483 56604
rect 7539 56602 7563 56604
rect 7619 56602 7643 56604
rect 7699 56602 7723 56604
rect 7779 56602 7785 56604
rect 7539 56550 7541 56602
rect 7721 56550 7723 56602
rect 7477 56548 7483 56550
rect 7539 56548 7563 56550
rect 7619 56548 7643 56550
rect 7699 56548 7723 56550
rect 7779 56548 7785 56550
rect 7477 56528 7785 56548
rect 7477 55516 7785 55536
rect 7477 55514 7483 55516
rect 7539 55514 7563 55516
rect 7619 55514 7643 55516
rect 7699 55514 7723 55516
rect 7779 55514 7785 55516
rect 7539 55462 7541 55514
rect 7721 55462 7723 55514
rect 7477 55460 7483 55462
rect 7539 55460 7563 55462
rect 7619 55460 7643 55462
rect 7699 55460 7723 55462
rect 7779 55460 7785 55462
rect 7477 55440 7785 55460
rect 7477 54428 7785 54448
rect 7477 54426 7483 54428
rect 7539 54426 7563 54428
rect 7619 54426 7643 54428
rect 7699 54426 7723 54428
rect 7779 54426 7785 54428
rect 7539 54374 7541 54426
rect 7721 54374 7723 54426
rect 7477 54372 7483 54374
rect 7539 54372 7563 54374
rect 7619 54372 7643 54374
rect 7699 54372 7723 54374
rect 7779 54372 7785 54374
rect 7477 54352 7785 54372
rect 7104 54120 7156 54126
rect 7104 54062 7156 54068
rect 7012 41676 7064 41682
rect 7012 41618 7064 41624
rect 6920 36848 6972 36854
rect 6920 36790 6972 36796
rect 7116 30802 7144 54062
rect 7477 53340 7785 53360
rect 7477 53338 7483 53340
rect 7539 53338 7563 53340
rect 7619 53338 7643 53340
rect 7699 53338 7723 53340
rect 7779 53338 7785 53340
rect 7539 53286 7541 53338
rect 7721 53286 7723 53338
rect 7477 53284 7483 53286
rect 7539 53284 7563 53286
rect 7619 53284 7643 53286
rect 7699 53284 7723 53286
rect 7779 53284 7785 53286
rect 7477 53264 7785 53284
rect 7288 53168 7340 53174
rect 7288 53110 7340 53116
rect 7196 50856 7248 50862
rect 7196 50798 7248 50804
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7208 11898 7236 50798
rect 7300 21894 7328 53110
rect 7380 53100 7432 53106
rect 7380 53042 7432 53048
rect 7392 23594 7420 53042
rect 7477 52252 7785 52272
rect 7477 52250 7483 52252
rect 7539 52250 7563 52252
rect 7619 52250 7643 52252
rect 7699 52250 7723 52252
rect 7779 52250 7785 52252
rect 7539 52198 7541 52250
rect 7721 52198 7723 52250
rect 7477 52196 7483 52198
rect 7539 52196 7563 52198
rect 7619 52196 7643 52198
rect 7699 52196 7723 52198
rect 7779 52196 7785 52198
rect 7477 52176 7785 52196
rect 7932 51468 7984 51474
rect 7932 51410 7984 51416
rect 7840 51332 7892 51338
rect 7840 51274 7892 51280
rect 7477 51164 7785 51184
rect 7477 51162 7483 51164
rect 7539 51162 7563 51164
rect 7619 51162 7643 51164
rect 7699 51162 7723 51164
rect 7779 51162 7785 51164
rect 7539 51110 7541 51162
rect 7721 51110 7723 51162
rect 7477 51108 7483 51110
rect 7539 51108 7563 51110
rect 7619 51108 7643 51110
rect 7699 51108 7723 51110
rect 7779 51108 7785 51110
rect 7477 51088 7785 51108
rect 7477 50076 7785 50096
rect 7477 50074 7483 50076
rect 7539 50074 7563 50076
rect 7619 50074 7643 50076
rect 7699 50074 7723 50076
rect 7779 50074 7785 50076
rect 7539 50022 7541 50074
rect 7721 50022 7723 50074
rect 7477 50020 7483 50022
rect 7539 50020 7563 50022
rect 7619 50020 7643 50022
rect 7699 50020 7723 50022
rect 7779 50020 7785 50022
rect 7477 50000 7785 50020
rect 7477 48988 7785 49008
rect 7477 48986 7483 48988
rect 7539 48986 7563 48988
rect 7619 48986 7643 48988
rect 7699 48986 7723 48988
rect 7779 48986 7785 48988
rect 7539 48934 7541 48986
rect 7721 48934 7723 48986
rect 7477 48932 7483 48934
rect 7539 48932 7563 48934
rect 7619 48932 7643 48934
rect 7699 48932 7723 48934
rect 7779 48932 7785 48934
rect 7477 48912 7785 48932
rect 7477 47900 7785 47920
rect 7477 47898 7483 47900
rect 7539 47898 7563 47900
rect 7619 47898 7643 47900
rect 7699 47898 7723 47900
rect 7779 47898 7785 47900
rect 7539 47846 7541 47898
rect 7721 47846 7723 47898
rect 7477 47844 7483 47846
rect 7539 47844 7563 47846
rect 7619 47844 7643 47846
rect 7699 47844 7723 47846
rect 7779 47844 7785 47846
rect 7477 47824 7785 47844
rect 7477 46812 7785 46832
rect 7477 46810 7483 46812
rect 7539 46810 7563 46812
rect 7619 46810 7643 46812
rect 7699 46810 7723 46812
rect 7779 46810 7785 46812
rect 7539 46758 7541 46810
rect 7721 46758 7723 46810
rect 7477 46756 7483 46758
rect 7539 46756 7563 46758
rect 7619 46756 7643 46758
rect 7699 46756 7723 46758
rect 7779 46756 7785 46758
rect 7477 46736 7785 46756
rect 7477 45724 7785 45744
rect 7477 45722 7483 45724
rect 7539 45722 7563 45724
rect 7619 45722 7643 45724
rect 7699 45722 7723 45724
rect 7779 45722 7785 45724
rect 7539 45670 7541 45722
rect 7721 45670 7723 45722
rect 7477 45668 7483 45670
rect 7539 45668 7563 45670
rect 7619 45668 7643 45670
rect 7699 45668 7723 45670
rect 7779 45668 7785 45670
rect 7477 45648 7785 45668
rect 7477 44636 7785 44656
rect 7477 44634 7483 44636
rect 7539 44634 7563 44636
rect 7619 44634 7643 44636
rect 7699 44634 7723 44636
rect 7779 44634 7785 44636
rect 7539 44582 7541 44634
rect 7721 44582 7723 44634
rect 7477 44580 7483 44582
rect 7539 44580 7563 44582
rect 7619 44580 7643 44582
rect 7699 44580 7723 44582
rect 7779 44580 7785 44582
rect 7477 44560 7785 44580
rect 7477 43548 7785 43568
rect 7477 43546 7483 43548
rect 7539 43546 7563 43548
rect 7619 43546 7643 43548
rect 7699 43546 7723 43548
rect 7779 43546 7785 43548
rect 7539 43494 7541 43546
rect 7721 43494 7723 43546
rect 7477 43492 7483 43494
rect 7539 43492 7563 43494
rect 7619 43492 7643 43494
rect 7699 43492 7723 43494
rect 7779 43492 7785 43494
rect 7477 43472 7785 43492
rect 7477 42460 7785 42480
rect 7477 42458 7483 42460
rect 7539 42458 7563 42460
rect 7619 42458 7643 42460
rect 7699 42458 7723 42460
rect 7779 42458 7785 42460
rect 7539 42406 7541 42458
rect 7721 42406 7723 42458
rect 7477 42404 7483 42406
rect 7539 42404 7563 42406
rect 7619 42404 7643 42406
rect 7699 42404 7723 42406
rect 7779 42404 7785 42406
rect 7477 42384 7785 42404
rect 7477 41372 7785 41392
rect 7477 41370 7483 41372
rect 7539 41370 7563 41372
rect 7619 41370 7643 41372
rect 7699 41370 7723 41372
rect 7779 41370 7785 41372
rect 7539 41318 7541 41370
rect 7721 41318 7723 41370
rect 7477 41316 7483 41318
rect 7539 41316 7563 41318
rect 7619 41316 7643 41318
rect 7699 41316 7723 41318
rect 7779 41316 7785 41318
rect 7477 41296 7785 41316
rect 7477 40284 7785 40304
rect 7477 40282 7483 40284
rect 7539 40282 7563 40284
rect 7619 40282 7643 40284
rect 7699 40282 7723 40284
rect 7779 40282 7785 40284
rect 7539 40230 7541 40282
rect 7721 40230 7723 40282
rect 7477 40228 7483 40230
rect 7539 40228 7563 40230
rect 7619 40228 7643 40230
rect 7699 40228 7723 40230
rect 7779 40228 7785 40230
rect 7477 40208 7785 40228
rect 7477 39196 7785 39216
rect 7477 39194 7483 39196
rect 7539 39194 7563 39196
rect 7619 39194 7643 39196
rect 7699 39194 7723 39196
rect 7779 39194 7785 39196
rect 7539 39142 7541 39194
rect 7721 39142 7723 39194
rect 7477 39140 7483 39142
rect 7539 39140 7563 39142
rect 7619 39140 7643 39142
rect 7699 39140 7723 39142
rect 7779 39140 7785 39142
rect 7477 39120 7785 39140
rect 7477 38108 7785 38128
rect 7477 38106 7483 38108
rect 7539 38106 7563 38108
rect 7619 38106 7643 38108
rect 7699 38106 7723 38108
rect 7779 38106 7785 38108
rect 7539 38054 7541 38106
rect 7721 38054 7723 38106
rect 7477 38052 7483 38054
rect 7539 38052 7563 38054
rect 7619 38052 7643 38054
rect 7699 38052 7723 38054
rect 7779 38052 7785 38054
rect 7477 38032 7785 38052
rect 7477 37020 7785 37040
rect 7477 37018 7483 37020
rect 7539 37018 7563 37020
rect 7619 37018 7643 37020
rect 7699 37018 7723 37020
rect 7779 37018 7785 37020
rect 7539 36966 7541 37018
rect 7721 36966 7723 37018
rect 7477 36964 7483 36966
rect 7539 36964 7563 36966
rect 7619 36964 7643 36966
rect 7699 36964 7723 36966
rect 7779 36964 7785 36966
rect 7477 36944 7785 36964
rect 7477 35932 7785 35952
rect 7477 35930 7483 35932
rect 7539 35930 7563 35932
rect 7619 35930 7643 35932
rect 7699 35930 7723 35932
rect 7779 35930 7785 35932
rect 7539 35878 7541 35930
rect 7721 35878 7723 35930
rect 7477 35876 7483 35878
rect 7539 35876 7563 35878
rect 7619 35876 7643 35878
rect 7699 35876 7723 35878
rect 7779 35876 7785 35878
rect 7477 35856 7785 35876
rect 7477 34844 7785 34864
rect 7477 34842 7483 34844
rect 7539 34842 7563 34844
rect 7619 34842 7643 34844
rect 7699 34842 7723 34844
rect 7779 34842 7785 34844
rect 7539 34790 7541 34842
rect 7721 34790 7723 34842
rect 7477 34788 7483 34790
rect 7539 34788 7563 34790
rect 7619 34788 7643 34790
rect 7699 34788 7723 34790
rect 7779 34788 7785 34790
rect 7477 34768 7785 34788
rect 7477 33756 7785 33776
rect 7477 33754 7483 33756
rect 7539 33754 7563 33756
rect 7619 33754 7643 33756
rect 7699 33754 7723 33756
rect 7779 33754 7785 33756
rect 7539 33702 7541 33754
rect 7721 33702 7723 33754
rect 7477 33700 7483 33702
rect 7539 33700 7563 33702
rect 7619 33700 7643 33702
rect 7699 33700 7723 33702
rect 7779 33700 7785 33702
rect 7477 33680 7785 33700
rect 7477 32668 7785 32688
rect 7477 32666 7483 32668
rect 7539 32666 7563 32668
rect 7619 32666 7643 32668
rect 7699 32666 7723 32668
rect 7779 32666 7785 32668
rect 7539 32614 7541 32666
rect 7721 32614 7723 32666
rect 7477 32612 7483 32614
rect 7539 32612 7563 32614
rect 7619 32612 7643 32614
rect 7699 32612 7723 32614
rect 7779 32612 7785 32614
rect 7477 32592 7785 32612
rect 7477 31580 7785 31600
rect 7477 31578 7483 31580
rect 7539 31578 7563 31580
rect 7619 31578 7643 31580
rect 7699 31578 7723 31580
rect 7779 31578 7785 31580
rect 7539 31526 7541 31578
rect 7721 31526 7723 31578
rect 7477 31524 7483 31526
rect 7539 31524 7563 31526
rect 7619 31524 7643 31526
rect 7699 31524 7723 31526
rect 7779 31524 7785 31526
rect 7477 31504 7785 31524
rect 7477 30492 7785 30512
rect 7477 30490 7483 30492
rect 7539 30490 7563 30492
rect 7619 30490 7643 30492
rect 7699 30490 7723 30492
rect 7779 30490 7785 30492
rect 7539 30438 7541 30490
rect 7721 30438 7723 30490
rect 7477 30436 7483 30438
rect 7539 30436 7563 30438
rect 7619 30436 7643 30438
rect 7699 30436 7723 30438
rect 7779 30436 7785 30438
rect 7477 30416 7785 30436
rect 7477 29404 7785 29424
rect 7477 29402 7483 29404
rect 7539 29402 7563 29404
rect 7619 29402 7643 29404
rect 7699 29402 7723 29404
rect 7779 29402 7785 29404
rect 7539 29350 7541 29402
rect 7721 29350 7723 29402
rect 7477 29348 7483 29350
rect 7539 29348 7563 29350
rect 7619 29348 7643 29350
rect 7699 29348 7723 29350
rect 7779 29348 7785 29350
rect 7477 29328 7785 29348
rect 7477 28316 7785 28336
rect 7477 28314 7483 28316
rect 7539 28314 7563 28316
rect 7619 28314 7643 28316
rect 7699 28314 7723 28316
rect 7779 28314 7785 28316
rect 7539 28262 7541 28314
rect 7721 28262 7723 28314
rect 7477 28260 7483 28262
rect 7539 28260 7563 28262
rect 7619 28260 7643 28262
rect 7699 28260 7723 28262
rect 7779 28260 7785 28262
rect 7477 28240 7785 28260
rect 7477 27228 7785 27248
rect 7477 27226 7483 27228
rect 7539 27226 7563 27228
rect 7619 27226 7643 27228
rect 7699 27226 7723 27228
rect 7779 27226 7785 27228
rect 7539 27174 7541 27226
rect 7721 27174 7723 27226
rect 7477 27172 7483 27174
rect 7539 27172 7563 27174
rect 7619 27172 7643 27174
rect 7699 27172 7723 27174
rect 7779 27172 7785 27174
rect 7477 27152 7785 27172
rect 7477 26140 7785 26160
rect 7477 26138 7483 26140
rect 7539 26138 7563 26140
rect 7619 26138 7643 26140
rect 7699 26138 7723 26140
rect 7779 26138 7785 26140
rect 7539 26086 7541 26138
rect 7721 26086 7723 26138
rect 7477 26084 7483 26086
rect 7539 26084 7563 26086
rect 7619 26084 7643 26086
rect 7699 26084 7723 26086
rect 7779 26084 7785 26086
rect 7477 26064 7785 26084
rect 7477 25052 7785 25072
rect 7477 25050 7483 25052
rect 7539 25050 7563 25052
rect 7619 25050 7643 25052
rect 7699 25050 7723 25052
rect 7779 25050 7785 25052
rect 7539 24998 7541 25050
rect 7721 24998 7723 25050
rect 7477 24996 7483 24998
rect 7539 24996 7563 24998
rect 7619 24996 7643 24998
rect 7699 24996 7723 24998
rect 7779 24996 7785 24998
rect 7477 24976 7785 24996
rect 7477 23964 7785 23984
rect 7477 23962 7483 23964
rect 7539 23962 7563 23964
rect 7619 23962 7643 23964
rect 7699 23962 7723 23964
rect 7779 23962 7785 23964
rect 7539 23910 7541 23962
rect 7721 23910 7723 23962
rect 7477 23908 7483 23910
rect 7539 23908 7563 23910
rect 7619 23908 7643 23910
rect 7699 23908 7723 23910
rect 7779 23908 7785 23910
rect 7477 23888 7785 23908
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7477 22876 7785 22896
rect 7477 22874 7483 22876
rect 7539 22874 7563 22876
rect 7619 22874 7643 22876
rect 7699 22874 7723 22876
rect 7779 22874 7785 22876
rect 7539 22822 7541 22874
rect 7721 22822 7723 22874
rect 7477 22820 7483 22822
rect 7539 22820 7563 22822
rect 7619 22820 7643 22822
rect 7699 22820 7723 22822
rect 7779 22820 7785 22822
rect 7477 22800 7785 22820
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 7477 21788 7785 21808
rect 7477 21786 7483 21788
rect 7539 21786 7563 21788
rect 7619 21786 7643 21788
rect 7699 21786 7723 21788
rect 7779 21786 7785 21788
rect 7539 21734 7541 21786
rect 7721 21734 7723 21786
rect 7477 21732 7483 21734
rect 7539 21732 7563 21734
rect 7619 21732 7643 21734
rect 7699 21732 7723 21734
rect 7779 21732 7785 21734
rect 7477 21712 7785 21732
rect 7477 20700 7785 20720
rect 7477 20698 7483 20700
rect 7539 20698 7563 20700
rect 7619 20698 7643 20700
rect 7699 20698 7723 20700
rect 7779 20698 7785 20700
rect 7539 20646 7541 20698
rect 7721 20646 7723 20698
rect 7477 20644 7483 20646
rect 7539 20644 7563 20646
rect 7619 20644 7643 20646
rect 7699 20644 7723 20646
rect 7779 20644 7785 20646
rect 7477 20624 7785 20644
rect 7477 19612 7785 19632
rect 7477 19610 7483 19612
rect 7539 19610 7563 19612
rect 7619 19610 7643 19612
rect 7699 19610 7723 19612
rect 7779 19610 7785 19612
rect 7539 19558 7541 19610
rect 7721 19558 7723 19610
rect 7477 19556 7483 19558
rect 7539 19556 7563 19558
rect 7619 19556 7643 19558
rect 7699 19556 7723 19558
rect 7779 19556 7785 19558
rect 7477 19536 7785 19556
rect 7477 18524 7785 18544
rect 7477 18522 7483 18524
rect 7539 18522 7563 18524
rect 7619 18522 7643 18524
rect 7699 18522 7723 18524
rect 7779 18522 7785 18524
rect 7539 18470 7541 18522
rect 7721 18470 7723 18522
rect 7477 18468 7483 18470
rect 7539 18468 7563 18470
rect 7619 18468 7643 18470
rect 7699 18468 7723 18470
rect 7779 18468 7785 18470
rect 7477 18448 7785 18468
rect 7477 17436 7785 17456
rect 7477 17434 7483 17436
rect 7539 17434 7563 17436
rect 7619 17434 7643 17436
rect 7699 17434 7723 17436
rect 7779 17434 7785 17436
rect 7539 17382 7541 17434
rect 7721 17382 7723 17434
rect 7477 17380 7483 17382
rect 7539 17380 7563 17382
rect 7619 17380 7643 17382
rect 7699 17380 7723 17382
rect 7779 17380 7785 17382
rect 7477 17360 7785 17380
rect 7477 16348 7785 16368
rect 7477 16346 7483 16348
rect 7539 16346 7563 16348
rect 7619 16346 7643 16348
rect 7699 16346 7723 16348
rect 7779 16346 7785 16348
rect 7539 16294 7541 16346
rect 7721 16294 7723 16346
rect 7477 16292 7483 16294
rect 7539 16292 7563 16294
rect 7619 16292 7643 16294
rect 7699 16292 7723 16294
rect 7779 16292 7785 16294
rect 7477 16272 7785 16292
rect 7477 15260 7785 15280
rect 7477 15258 7483 15260
rect 7539 15258 7563 15260
rect 7619 15258 7643 15260
rect 7699 15258 7723 15260
rect 7779 15258 7785 15260
rect 7539 15206 7541 15258
rect 7721 15206 7723 15258
rect 7477 15204 7483 15206
rect 7539 15204 7563 15206
rect 7619 15204 7643 15206
rect 7699 15204 7723 15206
rect 7779 15204 7785 15206
rect 7477 15184 7785 15204
rect 7477 14172 7785 14192
rect 7477 14170 7483 14172
rect 7539 14170 7563 14172
rect 7619 14170 7643 14172
rect 7699 14170 7723 14172
rect 7779 14170 7785 14172
rect 7539 14118 7541 14170
rect 7721 14118 7723 14170
rect 7477 14116 7483 14118
rect 7539 14116 7563 14118
rect 7619 14116 7643 14118
rect 7699 14116 7723 14118
rect 7779 14116 7785 14118
rect 7477 14096 7785 14116
rect 7477 13084 7785 13104
rect 7477 13082 7483 13084
rect 7539 13082 7563 13084
rect 7619 13082 7643 13084
rect 7699 13082 7723 13084
rect 7779 13082 7785 13084
rect 7539 13030 7541 13082
rect 7721 13030 7723 13082
rect 7477 13028 7483 13030
rect 7539 13028 7563 13030
rect 7619 13028 7643 13030
rect 7699 13028 7723 13030
rect 7779 13028 7785 13030
rect 7477 13008 7785 13028
rect 7852 12986 7880 51274
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12442 7972 51410
rect 8024 45960 8076 45966
rect 8024 45902 8076 45908
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7477 11996 7785 12016
rect 7477 11994 7483 11996
rect 7539 11994 7563 11996
rect 7619 11994 7643 11996
rect 7699 11994 7723 11996
rect 7779 11994 7785 11996
rect 7539 11942 7541 11994
rect 7721 11942 7723 11994
rect 7477 11940 7483 11942
rect 7539 11940 7563 11942
rect 7619 11940 7643 11942
rect 7699 11940 7723 11942
rect 7779 11940 7785 11942
rect 7477 11920 7785 11940
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7477 10908 7785 10928
rect 7477 10906 7483 10908
rect 7539 10906 7563 10908
rect 7619 10906 7643 10908
rect 7699 10906 7723 10908
rect 7779 10906 7785 10908
rect 7539 10854 7541 10906
rect 7721 10854 7723 10906
rect 7477 10852 7483 10854
rect 7539 10852 7563 10854
rect 7619 10852 7643 10854
rect 7699 10852 7723 10854
rect 7779 10852 7785 10854
rect 7477 10832 7785 10852
rect 7477 9820 7785 9840
rect 7477 9818 7483 9820
rect 7539 9818 7563 9820
rect 7619 9818 7643 9820
rect 7699 9818 7723 9820
rect 7779 9818 7785 9820
rect 7539 9766 7541 9818
rect 7721 9766 7723 9818
rect 7477 9764 7483 9766
rect 7539 9764 7563 9766
rect 7619 9764 7643 9766
rect 7699 9764 7723 9766
rect 7779 9764 7785 9766
rect 7477 9744 7785 9764
rect 7477 8732 7785 8752
rect 7477 8730 7483 8732
rect 7539 8730 7563 8732
rect 7619 8730 7643 8732
rect 7699 8730 7723 8732
rect 7779 8730 7785 8732
rect 7539 8678 7541 8730
rect 7721 8678 7723 8730
rect 7477 8676 7483 8678
rect 7539 8676 7563 8678
rect 7619 8676 7643 8678
rect 7699 8676 7723 8678
rect 7779 8676 7785 8678
rect 7477 8656 7785 8676
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 5845 8188 6153 8208
rect 5845 8186 5851 8188
rect 5907 8186 5931 8188
rect 5987 8186 6011 8188
rect 6067 8186 6091 8188
rect 6147 8186 6153 8188
rect 5907 8134 5909 8186
rect 6089 8134 6091 8186
rect 5845 8132 5851 8134
rect 5907 8132 5931 8134
rect 5987 8132 6011 8134
rect 6067 8132 6091 8134
rect 6147 8132 6153 8134
rect 5845 8112 6153 8132
rect 7477 7644 7785 7664
rect 7477 7642 7483 7644
rect 7539 7642 7563 7644
rect 7619 7642 7643 7644
rect 7699 7642 7723 7644
rect 7779 7642 7785 7644
rect 7539 7590 7541 7642
rect 7721 7590 7723 7642
rect 7477 7588 7483 7590
rect 7539 7588 7563 7590
rect 7619 7588 7643 7590
rect 7699 7588 7723 7590
rect 7779 7588 7785 7590
rect 7477 7568 7785 7588
rect 5845 7100 6153 7120
rect 5845 7098 5851 7100
rect 5907 7098 5931 7100
rect 5987 7098 6011 7100
rect 6067 7098 6091 7100
rect 6147 7098 6153 7100
rect 5907 7046 5909 7098
rect 6089 7046 6091 7098
rect 5845 7044 5851 7046
rect 5907 7044 5931 7046
rect 5987 7044 6011 7046
rect 6067 7044 6091 7046
rect 6147 7044 6153 7046
rect 5845 7024 6153 7044
rect 8036 6914 8064 45902
rect 8312 43722 8340 75414
rect 9968 75342 9996 76230
rect 10232 75880 10284 75886
rect 10232 75822 10284 75828
rect 10244 75721 10272 75822
rect 10230 75712 10286 75721
rect 10230 75647 10286 75656
rect 9956 75336 10008 75342
rect 9956 75278 10008 75284
rect 10140 75336 10192 75342
rect 10140 75278 10192 75284
rect 9956 75200 10008 75206
rect 9956 75142 10008 75148
rect 9968 74798 9996 75142
rect 10152 74905 10180 75278
rect 10138 74896 10194 74905
rect 10138 74831 10194 74840
rect 9956 74792 10008 74798
rect 9956 74734 10008 74740
rect 9109 74556 9417 74576
rect 9109 74554 9115 74556
rect 9171 74554 9195 74556
rect 9251 74554 9275 74556
rect 9331 74554 9355 74556
rect 9411 74554 9417 74556
rect 9171 74502 9173 74554
rect 9353 74502 9355 74554
rect 9109 74500 9115 74502
rect 9171 74500 9195 74502
rect 9251 74500 9275 74502
rect 9331 74500 9355 74502
rect 9411 74500 9417 74502
rect 9109 74480 9417 74500
rect 10140 74248 10192 74254
rect 10140 74190 10192 74196
rect 9956 74112 10008 74118
rect 10152 74089 10180 74190
rect 9956 74054 10008 74060
rect 10138 74080 10194 74089
rect 9864 73704 9916 73710
rect 9864 73646 9916 73652
rect 9109 73468 9417 73488
rect 9109 73466 9115 73468
rect 9171 73466 9195 73468
rect 9251 73466 9275 73468
rect 9331 73466 9355 73468
rect 9411 73466 9417 73468
rect 9171 73414 9173 73466
rect 9353 73414 9355 73466
rect 9109 73412 9115 73414
rect 9171 73412 9195 73414
rect 9251 73412 9275 73414
rect 9331 73412 9355 73414
rect 9411 73412 9417 73414
rect 9109 73392 9417 73412
rect 8392 72548 8444 72554
rect 8392 72490 8444 72496
rect 8300 43716 8352 43722
rect 8300 43658 8352 43664
rect 8404 41206 8432 72490
rect 9109 72380 9417 72400
rect 9109 72378 9115 72380
rect 9171 72378 9195 72380
rect 9251 72378 9275 72380
rect 9331 72378 9355 72380
rect 9411 72378 9417 72380
rect 9171 72326 9173 72378
rect 9353 72326 9355 72378
rect 9109 72324 9115 72326
rect 9171 72324 9195 72326
rect 9251 72324 9275 72326
rect 9331 72324 9355 72326
rect 9411 72324 9417 72326
rect 9109 72304 9417 72324
rect 9876 71738 9904 73646
rect 9968 72758 9996 74054
rect 10138 74015 10194 74024
rect 10140 73772 10192 73778
rect 10140 73714 10192 73720
rect 10152 73409 10180 73714
rect 10138 73400 10194 73409
rect 10138 73335 10194 73344
rect 9956 72752 10008 72758
rect 9956 72694 10008 72700
rect 10140 72684 10192 72690
rect 10140 72626 10192 72632
rect 9956 72616 10008 72622
rect 10152 72593 10180 72626
rect 9956 72558 10008 72564
rect 10138 72584 10194 72593
rect 9968 72282 9996 72558
rect 10138 72519 10194 72528
rect 9956 72276 10008 72282
rect 9956 72218 10008 72224
rect 10140 72072 10192 72078
rect 10140 72014 10192 72020
rect 10152 71777 10180 72014
rect 10138 71768 10194 71777
rect 9864 71732 9916 71738
rect 10138 71703 10194 71712
rect 9864 71674 9916 71680
rect 10140 71596 10192 71602
rect 10140 71538 10192 71544
rect 9109 71292 9417 71312
rect 9109 71290 9115 71292
rect 9171 71290 9195 71292
rect 9251 71290 9275 71292
rect 9331 71290 9355 71292
rect 9411 71290 9417 71292
rect 9171 71238 9173 71290
rect 9353 71238 9355 71290
rect 9109 71236 9115 71238
rect 9171 71236 9195 71238
rect 9251 71236 9275 71238
rect 9331 71236 9355 71238
rect 9411 71236 9417 71238
rect 9109 71216 9417 71236
rect 10152 71097 10180 71538
rect 10138 71088 10194 71097
rect 10138 71023 10194 71032
rect 10140 70372 10192 70378
rect 10140 70314 10192 70320
rect 10152 70281 10180 70314
rect 10138 70272 10194 70281
rect 9109 70204 9417 70224
rect 10138 70207 10194 70216
rect 9109 70202 9115 70204
rect 9171 70202 9195 70204
rect 9251 70202 9275 70204
rect 9331 70202 9355 70204
rect 9411 70202 9417 70204
rect 9171 70150 9173 70202
rect 9353 70150 9355 70202
rect 9109 70148 9115 70150
rect 9171 70148 9195 70150
rect 9251 70148 9275 70150
rect 9331 70148 9355 70150
rect 9411 70148 9417 70150
rect 9109 70128 9417 70148
rect 10140 69896 10192 69902
rect 10140 69838 10192 69844
rect 10152 69465 10180 69838
rect 10138 69456 10194 69465
rect 10138 69391 10194 69400
rect 9956 69352 10008 69358
rect 9956 69294 10008 69300
rect 9109 69116 9417 69136
rect 9109 69114 9115 69116
rect 9171 69114 9195 69116
rect 9251 69114 9275 69116
rect 9331 69114 9355 69116
rect 9411 69114 9417 69116
rect 9171 69062 9173 69114
rect 9353 69062 9355 69114
rect 9109 69060 9115 69062
rect 9171 69060 9195 69062
rect 9251 69060 9275 69062
rect 9331 69060 9355 69062
rect 9411 69060 9417 69062
rect 9109 69040 9417 69060
rect 9968 69018 9996 69294
rect 9956 69012 10008 69018
rect 9956 68954 10008 68960
rect 10140 68808 10192 68814
rect 10138 68776 10140 68785
rect 10192 68776 10194 68785
rect 10138 68711 10194 68720
rect 10140 68332 10192 68338
rect 10140 68274 10192 68280
rect 9109 68028 9417 68048
rect 9109 68026 9115 68028
rect 9171 68026 9195 68028
rect 9251 68026 9275 68028
rect 9331 68026 9355 68028
rect 9411 68026 9417 68028
rect 9171 67974 9173 68026
rect 9353 67974 9355 68026
rect 9109 67972 9115 67974
rect 9171 67972 9195 67974
rect 9251 67972 9275 67974
rect 9331 67972 9355 67974
rect 9411 67972 9417 67974
rect 9109 67952 9417 67972
rect 10152 67969 10180 68274
rect 10138 67960 10194 67969
rect 10138 67895 10194 67904
rect 10140 67244 10192 67250
rect 10140 67186 10192 67192
rect 10152 67153 10180 67186
rect 10138 67144 10194 67153
rect 10138 67079 10194 67088
rect 9956 67040 10008 67046
rect 9956 66982 10008 66988
rect 9109 66940 9417 66960
rect 9109 66938 9115 66940
rect 9171 66938 9195 66940
rect 9251 66938 9275 66940
rect 9331 66938 9355 66940
rect 9411 66938 9417 66940
rect 9171 66886 9173 66938
rect 9353 66886 9355 66938
rect 9109 66884 9115 66886
rect 9171 66884 9195 66886
rect 9251 66884 9275 66886
rect 9331 66884 9355 66886
rect 9411 66884 9417 66886
rect 9109 66864 9417 66884
rect 9864 66496 9916 66502
rect 9864 66438 9916 66444
rect 9109 65852 9417 65872
rect 9109 65850 9115 65852
rect 9171 65850 9195 65852
rect 9251 65850 9275 65852
rect 9331 65850 9355 65852
rect 9411 65850 9417 65852
rect 9171 65798 9173 65850
rect 9353 65798 9355 65850
rect 9109 65796 9115 65798
rect 9171 65796 9195 65798
rect 9251 65796 9275 65798
rect 9331 65796 9355 65798
rect 9411 65796 9417 65798
rect 9109 65776 9417 65796
rect 9876 65618 9904 66438
rect 9968 66230 9996 66982
rect 10140 66632 10192 66638
rect 10140 66574 10192 66580
rect 10152 66473 10180 66574
rect 10138 66464 10194 66473
rect 10138 66399 10194 66408
rect 9956 66224 10008 66230
rect 9956 66166 10008 66172
rect 10140 66156 10192 66162
rect 10140 66098 10192 66104
rect 10152 65657 10180 66098
rect 10138 65648 10194 65657
rect 9864 65612 9916 65618
rect 10138 65583 10194 65592
rect 9864 65554 9916 65560
rect 10140 65068 10192 65074
rect 10140 65010 10192 65016
rect 10152 64841 10180 65010
rect 10138 64832 10194 64841
rect 9109 64764 9417 64784
rect 10138 64767 10194 64776
rect 9109 64762 9115 64764
rect 9171 64762 9195 64764
rect 9251 64762 9275 64764
rect 9331 64762 9355 64764
rect 9411 64762 9417 64764
rect 9171 64710 9173 64762
rect 9353 64710 9355 64762
rect 9109 64708 9115 64710
rect 9171 64708 9195 64710
rect 9251 64708 9275 64710
rect 9331 64708 9355 64710
rect 9411 64708 9417 64710
rect 9109 64688 9417 64708
rect 10140 64456 10192 64462
rect 10140 64398 10192 64404
rect 9956 64320 10008 64326
rect 9956 64262 10008 64268
rect 9109 63676 9417 63696
rect 9109 63674 9115 63676
rect 9171 63674 9195 63676
rect 9251 63674 9275 63676
rect 9331 63674 9355 63676
rect 9411 63674 9417 63676
rect 9171 63622 9173 63674
rect 9353 63622 9355 63674
rect 9109 63620 9115 63622
rect 9171 63620 9195 63622
rect 9251 63620 9275 63622
rect 9331 63620 9355 63622
rect 9411 63620 9417 63622
rect 9109 63600 9417 63620
rect 9864 63232 9916 63238
rect 9864 63174 9916 63180
rect 8484 62756 8536 62762
rect 8484 62698 8536 62704
rect 8392 41200 8444 41206
rect 8392 41142 8444 41148
rect 8496 36718 8524 62698
rect 9109 62588 9417 62608
rect 9109 62586 9115 62588
rect 9171 62586 9195 62588
rect 9251 62586 9275 62588
rect 9331 62586 9355 62588
rect 9411 62586 9417 62588
rect 9171 62534 9173 62586
rect 9353 62534 9355 62586
rect 9109 62532 9115 62534
rect 9171 62532 9195 62534
rect 9251 62532 9275 62534
rect 9331 62532 9355 62534
rect 9411 62532 9417 62534
rect 9109 62512 9417 62532
rect 9772 62144 9824 62150
rect 9772 62086 9824 62092
rect 9109 61500 9417 61520
rect 9109 61498 9115 61500
rect 9171 61498 9195 61500
rect 9251 61498 9275 61500
rect 9331 61498 9355 61500
rect 9411 61498 9417 61500
rect 9171 61446 9173 61498
rect 9353 61446 9355 61498
rect 9109 61444 9115 61446
rect 9171 61444 9195 61446
rect 9251 61444 9275 61446
rect 9331 61444 9355 61446
rect 9411 61444 9417 61446
rect 9109 61424 9417 61444
rect 9109 60412 9417 60432
rect 9109 60410 9115 60412
rect 9171 60410 9195 60412
rect 9251 60410 9275 60412
rect 9331 60410 9355 60412
rect 9411 60410 9417 60412
rect 9171 60358 9173 60410
rect 9353 60358 9355 60410
rect 9109 60356 9115 60358
rect 9171 60356 9195 60358
rect 9251 60356 9275 60358
rect 9331 60356 9355 60358
rect 9411 60356 9417 60358
rect 9109 60336 9417 60356
rect 9784 59702 9812 62086
rect 9876 60790 9904 63174
rect 9968 62966 9996 64262
rect 10152 64161 10180 64398
rect 10138 64152 10194 64161
rect 10138 64087 10194 64096
rect 10140 63368 10192 63374
rect 10138 63336 10140 63345
rect 10192 63336 10194 63345
rect 10138 63271 10194 63280
rect 9956 62960 10008 62966
rect 9956 62902 10008 62908
rect 10140 62892 10192 62898
rect 10140 62834 10192 62840
rect 10152 62529 10180 62834
rect 10138 62520 10194 62529
rect 10138 62455 10194 62464
rect 10140 62280 10192 62286
rect 10140 62222 10192 62228
rect 10152 61849 10180 62222
rect 10138 61840 10194 61849
rect 10138 61775 10194 61784
rect 10140 61192 10192 61198
rect 10140 61134 10192 61140
rect 9956 61056 10008 61062
rect 10152 61033 10180 61134
rect 9956 60998 10008 61004
rect 10138 61024 10194 61033
rect 9864 60784 9916 60790
rect 9864 60726 9916 60732
rect 9968 60602 9996 60998
rect 10138 60959 10194 60968
rect 10140 60716 10192 60722
rect 10140 60658 10192 60664
rect 9876 60574 9996 60602
rect 9876 60042 9904 60574
rect 9956 60512 10008 60518
rect 9956 60454 10008 60460
rect 9864 60036 9916 60042
rect 9864 59978 9916 59984
rect 9772 59696 9824 59702
rect 9772 59638 9824 59644
rect 9109 59324 9417 59344
rect 9109 59322 9115 59324
rect 9171 59322 9195 59324
rect 9251 59322 9275 59324
rect 9331 59322 9355 59324
rect 9411 59322 9417 59324
rect 9171 59270 9173 59322
rect 9353 59270 9355 59322
rect 9109 59268 9115 59270
rect 9171 59268 9195 59270
rect 9251 59268 9275 59270
rect 9331 59268 9355 59270
rect 9411 59268 9417 59270
rect 9109 59248 9417 59268
rect 9968 59022 9996 60454
rect 10152 60353 10180 60658
rect 10138 60344 10194 60353
rect 10138 60279 10194 60288
rect 10140 59628 10192 59634
rect 10140 59570 10192 59576
rect 10152 59537 10180 59570
rect 10138 59528 10194 59537
rect 10138 59463 10194 59472
rect 9956 59016 10008 59022
rect 9956 58958 10008 58964
rect 10140 59016 10192 59022
rect 10140 58958 10192 58964
rect 9956 58880 10008 58886
rect 9956 58822 10008 58828
rect 8576 58404 8628 58410
rect 8576 58346 8628 58352
rect 8484 36712 8536 36718
rect 8484 36654 8536 36660
rect 8588 34134 8616 58346
rect 9109 58236 9417 58256
rect 9109 58234 9115 58236
rect 9171 58234 9195 58236
rect 9251 58234 9275 58236
rect 9331 58234 9355 58236
rect 9411 58234 9417 58236
rect 9171 58182 9173 58234
rect 9353 58182 9355 58234
rect 9109 58180 9115 58182
rect 9171 58180 9195 58182
rect 9251 58180 9275 58182
rect 9331 58180 9355 58182
rect 9411 58180 9417 58182
rect 9109 58160 9417 58180
rect 9968 57866 9996 58822
rect 10152 58721 10180 58958
rect 10138 58712 10194 58721
rect 10138 58647 10194 58656
rect 10140 58472 10192 58478
rect 10140 58414 10192 58420
rect 10152 58041 10180 58414
rect 10138 58032 10194 58041
rect 10138 57967 10194 57976
rect 9956 57860 10008 57866
rect 9956 57802 10008 57808
rect 10140 57384 10192 57390
rect 10140 57326 10192 57332
rect 10152 57225 10180 57326
rect 10138 57216 10194 57225
rect 9109 57148 9417 57168
rect 10138 57151 10194 57160
rect 9109 57146 9115 57148
rect 9171 57146 9195 57148
rect 9251 57146 9275 57148
rect 9331 57146 9355 57148
rect 9411 57146 9417 57148
rect 9171 57094 9173 57146
rect 9353 57094 9355 57146
rect 9109 57092 9115 57094
rect 9171 57092 9195 57094
rect 9251 57092 9275 57094
rect 9331 57092 9355 57094
rect 9411 57092 9417 57094
rect 9109 57072 9417 57092
rect 10140 56840 10192 56846
rect 10140 56782 10192 56788
rect 8852 56500 8904 56506
rect 8852 56442 8904 56448
rect 8760 55820 8812 55826
rect 8760 55762 8812 55768
rect 8668 53712 8720 53718
rect 8668 53654 8720 53660
rect 8576 34128 8628 34134
rect 8576 34070 8628 34076
rect 8680 30870 8708 53654
rect 8772 34678 8800 55762
rect 8864 35222 8892 56442
rect 10152 56409 10180 56782
rect 10138 56400 10194 56409
rect 10138 56335 10194 56344
rect 9864 56160 9916 56166
rect 9864 56102 9916 56108
rect 9109 56060 9417 56080
rect 9109 56058 9115 56060
rect 9171 56058 9195 56060
rect 9251 56058 9275 56060
rect 9331 56058 9355 56060
rect 9411 56058 9417 56060
rect 9171 56006 9173 56058
rect 9353 56006 9355 56058
rect 9109 56004 9115 56006
rect 9171 56004 9195 56006
rect 9251 56004 9275 56006
rect 9331 56004 9355 56006
rect 9411 56004 9417 56006
rect 9109 55984 9417 56004
rect 9109 54972 9417 54992
rect 9109 54970 9115 54972
rect 9171 54970 9195 54972
rect 9251 54970 9275 54972
rect 9331 54970 9355 54972
rect 9411 54970 9417 54972
rect 9171 54918 9173 54970
rect 9353 54918 9355 54970
rect 9109 54916 9115 54918
rect 9171 54916 9195 54918
rect 9251 54916 9275 54918
rect 9331 54916 9355 54918
rect 9411 54916 9417 54918
rect 9109 54896 9417 54916
rect 9876 54194 9904 56102
rect 10140 55752 10192 55758
rect 10138 55720 10140 55729
rect 10192 55720 10194 55729
rect 10138 55655 10194 55664
rect 10232 55208 10284 55214
rect 10232 55150 10284 55156
rect 9956 55072 10008 55078
rect 9956 55014 10008 55020
rect 9864 54188 9916 54194
rect 9864 54130 9916 54136
rect 9864 53984 9916 53990
rect 9864 53926 9916 53932
rect 9109 53884 9417 53904
rect 9109 53882 9115 53884
rect 9171 53882 9195 53884
rect 9251 53882 9275 53884
rect 9331 53882 9355 53884
rect 9411 53882 9417 53884
rect 9171 53830 9173 53882
rect 9353 53830 9355 53882
rect 9109 53828 9115 53830
rect 9171 53828 9195 53830
rect 9251 53828 9275 53830
rect 9331 53828 9355 53830
rect 9411 53828 9417 53830
rect 9109 53808 9417 53828
rect 9876 53106 9904 53926
rect 9968 53514 9996 55014
rect 10244 54913 10272 55150
rect 10230 54904 10286 54913
rect 10230 54839 10286 54848
rect 10046 54088 10102 54097
rect 10046 54023 10048 54032
rect 10100 54023 10102 54032
rect 10048 53994 10100 54000
rect 9956 53508 10008 53514
rect 9956 53450 10008 53456
rect 10048 53440 10100 53446
rect 10046 53408 10048 53417
rect 10100 53408 10102 53417
rect 10046 53343 10102 53352
rect 9864 53100 9916 53106
rect 9864 53042 9916 53048
rect 10048 52896 10100 52902
rect 10048 52838 10100 52844
rect 9109 52796 9417 52816
rect 9109 52794 9115 52796
rect 9171 52794 9195 52796
rect 9251 52794 9275 52796
rect 9331 52794 9355 52796
rect 9411 52794 9417 52796
rect 9171 52742 9173 52794
rect 9353 52742 9355 52794
rect 9109 52740 9115 52742
rect 9171 52740 9195 52742
rect 9251 52740 9275 52742
rect 9331 52740 9355 52742
rect 9411 52740 9417 52742
rect 9109 52720 9417 52740
rect 10060 52601 10088 52838
rect 10046 52592 10102 52601
rect 10046 52527 10102 52536
rect 10048 51808 10100 51814
rect 10046 51776 10048 51785
rect 10100 51776 10102 51785
rect 9109 51708 9417 51728
rect 10046 51711 10102 51720
rect 9109 51706 9115 51708
rect 9171 51706 9195 51708
rect 9251 51706 9275 51708
rect 9331 51706 9355 51708
rect 9411 51706 9417 51708
rect 9171 51654 9173 51706
rect 9353 51654 9355 51706
rect 9109 51652 9115 51654
rect 9171 51652 9195 51654
rect 9251 51652 9275 51654
rect 9331 51652 9355 51654
rect 9411 51652 9417 51654
rect 9109 51632 9417 51652
rect 9864 51400 9916 51406
rect 9864 51342 9916 51348
rect 9876 51066 9904 51342
rect 10048 51264 10100 51270
rect 10048 51206 10100 51212
rect 10060 51105 10088 51206
rect 10046 51096 10102 51105
rect 9864 51060 9916 51066
rect 10046 51031 10102 51040
rect 9864 51002 9916 51008
rect 9109 50620 9417 50640
rect 9109 50618 9115 50620
rect 9171 50618 9195 50620
rect 9251 50618 9275 50620
rect 9331 50618 9355 50620
rect 9411 50618 9417 50620
rect 9171 50566 9173 50618
rect 9353 50566 9355 50618
rect 9109 50564 9115 50566
rect 9171 50564 9195 50566
rect 9251 50564 9275 50566
rect 9331 50564 9355 50566
rect 9411 50564 9417 50566
rect 9109 50544 9417 50564
rect 10046 50280 10102 50289
rect 10046 50215 10102 50224
rect 10060 50182 10088 50215
rect 10048 50176 10100 50182
rect 10048 50118 10100 50124
rect 9864 49836 9916 49842
rect 9864 49778 9916 49784
rect 9109 49532 9417 49552
rect 9109 49530 9115 49532
rect 9171 49530 9195 49532
rect 9251 49530 9275 49532
rect 9331 49530 9355 49532
rect 9411 49530 9417 49532
rect 9171 49478 9173 49530
rect 9353 49478 9355 49530
rect 9109 49476 9115 49478
rect 9171 49476 9195 49478
rect 9251 49476 9275 49478
rect 9331 49476 9355 49478
rect 9411 49476 9417 49478
rect 9109 49456 9417 49476
rect 9772 49224 9824 49230
rect 9772 49166 9824 49172
rect 9109 48444 9417 48464
rect 9109 48442 9115 48444
rect 9171 48442 9195 48444
rect 9251 48442 9275 48444
rect 9331 48442 9355 48444
rect 9411 48442 9417 48444
rect 9171 48390 9173 48442
rect 9353 48390 9355 48442
rect 9109 48388 9115 48390
rect 9171 48388 9195 48390
rect 9251 48388 9275 48390
rect 9331 48388 9355 48390
rect 9411 48388 9417 48390
rect 9109 48368 9417 48388
rect 9109 47356 9417 47376
rect 9109 47354 9115 47356
rect 9171 47354 9195 47356
rect 9251 47354 9275 47356
rect 9331 47354 9355 47356
rect 9411 47354 9417 47356
rect 9171 47302 9173 47354
rect 9353 47302 9355 47354
rect 9109 47300 9115 47302
rect 9171 47300 9195 47302
rect 9251 47300 9275 47302
rect 9331 47300 9355 47302
rect 9411 47300 9417 47302
rect 9109 47280 9417 47300
rect 8944 46640 8996 46646
rect 8944 46582 8996 46588
rect 8852 35216 8904 35222
rect 8852 35158 8904 35164
rect 8760 34672 8812 34678
rect 8760 34614 8812 34620
rect 8668 30864 8720 30870
rect 8668 30806 8720 30812
rect 8956 23526 8984 46582
rect 9036 46504 9088 46510
rect 9036 46446 9088 46452
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 9048 10742 9076 46446
rect 9784 46442 9812 49166
rect 9876 48006 9904 49778
rect 10048 49632 10100 49638
rect 10048 49574 10100 49580
rect 10060 49473 10088 49574
rect 10046 49464 10102 49473
rect 10046 49399 10102 49408
rect 10048 49088 10100 49094
rect 10048 49030 10100 49036
rect 10060 48793 10088 49030
rect 10046 48784 10102 48793
rect 10046 48719 10102 48728
rect 9864 48000 9916 48006
rect 10048 48000 10100 48006
rect 9864 47942 9916 47948
rect 10046 47968 10048 47977
rect 10100 47968 10102 47977
rect 10046 47903 10102 47912
rect 10048 47456 10100 47462
rect 10048 47398 10100 47404
rect 10060 47161 10088 47398
rect 10046 47152 10102 47161
rect 10046 47087 10102 47096
rect 10046 46472 10102 46481
rect 9772 46436 9824 46442
rect 10046 46407 10048 46416
rect 9772 46378 9824 46384
rect 10100 46407 10102 46416
rect 10048 46378 10100 46384
rect 9109 46268 9417 46288
rect 9109 46266 9115 46268
rect 9171 46266 9195 46268
rect 9251 46266 9275 46268
rect 9331 46266 9355 46268
rect 9411 46266 9417 46268
rect 9171 46214 9173 46266
rect 9353 46214 9355 46266
rect 9109 46212 9115 46214
rect 9171 46212 9195 46214
rect 9251 46212 9275 46214
rect 9331 46212 9355 46214
rect 9411 46212 9417 46214
rect 9109 46192 9417 46212
rect 9864 45960 9916 45966
rect 9864 45902 9916 45908
rect 9109 45180 9417 45200
rect 9109 45178 9115 45180
rect 9171 45178 9195 45180
rect 9251 45178 9275 45180
rect 9331 45178 9355 45180
rect 9411 45178 9417 45180
rect 9171 45126 9173 45178
rect 9353 45126 9355 45178
rect 9109 45124 9115 45126
rect 9171 45124 9195 45126
rect 9251 45124 9275 45126
rect 9331 45124 9355 45126
rect 9411 45124 9417 45126
rect 9109 45104 9417 45124
rect 9680 44872 9732 44878
rect 9680 44814 9732 44820
rect 9692 44334 9720 44814
rect 9772 44396 9824 44402
rect 9772 44338 9824 44344
rect 9680 44328 9732 44334
rect 9680 44270 9732 44276
rect 9109 44092 9417 44112
rect 9109 44090 9115 44092
rect 9171 44090 9195 44092
rect 9251 44090 9275 44092
rect 9331 44090 9355 44092
rect 9411 44090 9417 44092
rect 9171 44038 9173 44090
rect 9353 44038 9355 44090
rect 9109 44036 9115 44038
rect 9171 44036 9195 44038
rect 9251 44036 9275 44038
rect 9331 44036 9355 44038
rect 9411 44036 9417 44038
rect 9109 44016 9417 44036
rect 9588 43784 9640 43790
rect 9588 43726 9640 43732
rect 9109 43004 9417 43024
rect 9109 43002 9115 43004
rect 9171 43002 9195 43004
rect 9251 43002 9275 43004
rect 9331 43002 9355 43004
rect 9411 43002 9417 43004
rect 9171 42950 9173 43002
rect 9353 42950 9355 43002
rect 9109 42948 9115 42950
rect 9171 42948 9195 42950
rect 9251 42948 9275 42950
rect 9331 42948 9355 42950
rect 9411 42948 9417 42950
rect 9109 42928 9417 42948
rect 9600 42362 9628 43726
rect 9680 43648 9732 43654
rect 9680 43590 9732 43596
rect 9692 42838 9720 43590
rect 9784 43382 9812 44338
rect 9876 43450 9904 45902
rect 10048 45824 10100 45830
rect 10048 45766 10100 45772
rect 10060 45665 10088 45766
rect 10046 45656 10102 45665
rect 10046 45591 10102 45600
rect 10046 44840 10102 44849
rect 10046 44775 10102 44784
rect 10060 44742 10088 44775
rect 10048 44736 10100 44742
rect 10048 44678 10100 44684
rect 10048 44192 10100 44198
rect 10046 44160 10048 44169
rect 10100 44160 10102 44169
rect 10046 44095 10102 44104
rect 10048 43648 10100 43654
rect 10048 43590 10100 43596
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9772 43376 9824 43382
rect 10060 43353 10088 43590
rect 9772 43318 9824 43324
rect 10046 43344 10102 43353
rect 10046 43279 10102 43288
rect 9680 42832 9732 42838
rect 9680 42774 9732 42780
rect 10048 42560 10100 42566
rect 10046 42528 10048 42537
rect 10100 42528 10102 42537
rect 10046 42463 10102 42472
rect 9588 42356 9640 42362
rect 9588 42298 9640 42304
rect 9864 42220 9916 42226
rect 9864 42162 9916 42168
rect 9109 41916 9417 41936
rect 9109 41914 9115 41916
rect 9171 41914 9195 41916
rect 9251 41914 9275 41916
rect 9331 41914 9355 41916
rect 9411 41914 9417 41916
rect 9171 41862 9173 41914
rect 9353 41862 9355 41914
rect 9109 41860 9115 41862
rect 9171 41860 9195 41862
rect 9251 41860 9275 41862
rect 9331 41860 9355 41862
rect 9411 41860 9417 41862
rect 9109 41840 9417 41860
rect 9876 41818 9904 42162
rect 10048 42016 10100 42022
rect 10048 41958 10100 41964
rect 10060 41857 10088 41958
rect 10046 41848 10102 41857
rect 9864 41812 9916 41818
rect 10046 41783 10102 41792
rect 9864 41754 9916 41760
rect 9680 41132 9732 41138
rect 9680 41074 9732 41080
rect 9109 40828 9417 40848
rect 9109 40826 9115 40828
rect 9171 40826 9195 40828
rect 9251 40826 9275 40828
rect 9331 40826 9355 40828
rect 9411 40826 9417 40828
rect 9171 40774 9173 40826
rect 9353 40774 9355 40826
rect 9109 40772 9115 40774
rect 9171 40772 9195 40774
rect 9251 40772 9275 40774
rect 9331 40772 9355 40774
rect 9411 40772 9417 40774
rect 9109 40752 9417 40772
rect 9692 39914 9720 41074
rect 10046 41032 10102 41041
rect 10046 40967 10048 40976
rect 10100 40967 10102 40976
rect 10048 40938 10100 40944
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 9772 40044 9824 40050
rect 9772 39986 9824 39992
rect 9680 39908 9732 39914
rect 9680 39850 9732 39856
rect 9109 39740 9417 39760
rect 9109 39738 9115 39740
rect 9171 39738 9195 39740
rect 9251 39738 9275 39740
rect 9331 39738 9355 39740
rect 9411 39738 9417 39740
rect 9171 39686 9173 39738
rect 9353 39686 9355 39738
rect 9109 39684 9115 39686
rect 9171 39684 9195 39686
rect 9251 39684 9275 39686
rect 9331 39684 9355 39686
rect 9411 39684 9417 39686
rect 9109 39664 9417 39684
rect 9109 38652 9417 38672
rect 9109 38650 9115 38652
rect 9171 38650 9195 38652
rect 9251 38650 9275 38652
rect 9331 38650 9355 38652
rect 9411 38650 9417 38652
rect 9171 38598 9173 38650
rect 9353 38598 9355 38650
rect 9109 38596 9115 38598
rect 9171 38596 9195 38598
rect 9251 38596 9275 38598
rect 9331 38596 9355 38598
rect 9411 38596 9417 38598
rect 9109 38576 9417 38596
rect 9784 38554 9812 39986
rect 9876 39098 9904 40462
rect 10048 40384 10100 40390
rect 10046 40352 10048 40361
rect 10100 40352 10102 40361
rect 10046 40287 10102 40296
rect 10048 39840 10100 39846
rect 10048 39782 10100 39788
rect 10060 39545 10088 39782
rect 10046 39536 10102 39545
rect 10046 39471 10102 39480
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 9864 38956 9916 38962
rect 9864 38898 9916 38904
rect 9772 38548 9824 38554
rect 9772 38490 9824 38496
rect 9109 37564 9417 37584
rect 9109 37562 9115 37564
rect 9171 37562 9195 37564
rect 9251 37562 9275 37564
rect 9331 37562 9355 37564
rect 9411 37562 9417 37564
rect 9171 37510 9173 37562
rect 9353 37510 9355 37562
rect 9109 37508 9115 37510
rect 9171 37508 9195 37510
rect 9251 37508 9275 37510
rect 9331 37508 9355 37510
rect 9411 37508 9417 37510
rect 9109 37488 9417 37508
rect 9876 37398 9904 38898
rect 10048 38752 10100 38758
rect 10046 38720 10048 38729
rect 10100 38720 10102 38729
rect 10046 38655 10102 38664
rect 10048 38208 10100 38214
rect 10048 38150 10100 38156
rect 10060 38049 10088 38150
rect 10046 38040 10102 38049
rect 10046 37975 10102 37984
rect 9864 37392 9916 37398
rect 9864 37334 9916 37340
rect 10046 37224 10102 37233
rect 10046 37159 10102 37168
rect 10060 37126 10088 37159
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 9772 36780 9824 36786
rect 9772 36722 9824 36728
rect 9109 36476 9417 36496
rect 9109 36474 9115 36476
rect 9171 36474 9195 36476
rect 9251 36474 9275 36476
rect 9331 36474 9355 36476
rect 9411 36474 9417 36476
rect 9171 36422 9173 36474
rect 9353 36422 9355 36474
rect 9109 36420 9115 36422
rect 9171 36420 9195 36422
rect 9251 36420 9275 36422
rect 9331 36420 9355 36422
rect 9411 36420 9417 36422
rect 9109 36400 9417 36420
rect 9109 35388 9417 35408
rect 9109 35386 9115 35388
rect 9171 35386 9195 35388
rect 9251 35386 9275 35388
rect 9331 35386 9355 35388
rect 9411 35386 9417 35388
rect 9171 35334 9173 35386
rect 9353 35334 9355 35386
rect 9109 35332 9115 35334
rect 9171 35332 9195 35334
rect 9251 35332 9275 35334
rect 9331 35332 9355 35334
rect 9411 35332 9417 35334
rect 9109 35312 9417 35332
rect 9680 34604 9732 34610
rect 9680 34546 9732 34552
rect 9109 34300 9417 34320
rect 9109 34298 9115 34300
rect 9171 34298 9195 34300
rect 9251 34298 9275 34300
rect 9331 34298 9355 34300
rect 9411 34298 9417 34300
rect 9171 34246 9173 34298
rect 9353 34246 9355 34298
rect 9109 34244 9115 34246
rect 9171 34244 9195 34246
rect 9251 34244 9275 34246
rect 9331 34244 9355 34246
rect 9411 34244 9417 34246
rect 9109 34224 9417 34244
rect 9109 33212 9417 33232
rect 9109 33210 9115 33212
rect 9171 33210 9195 33212
rect 9251 33210 9275 33212
rect 9331 33210 9355 33212
rect 9411 33210 9417 33212
rect 9171 33158 9173 33210
rect 9353 33158 9355 33210
rect 9109 33156 9115 33158
rect 9171 33156 9195 33158
rect 9251 33156 9275 33158
rect 9331 33156 9355 33158
rect 9411 33156 9417 33158
rect 9109 33136 9417 33156
rect 9692 33046 9720 34546
rect 9784 34202 9812 36722
rect 10048 36576 10100 36582
rect 10048 36518 10100 36524
rect 10060 36417 10088 36518
rect 10046 36408 10102 36417
rect 10046 36343 10102 36352
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 9876 35290 9904 36110
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 10060 35737 10088 35974
rect 10046 35728 10102 35737
rect 10046 35663 10102 35672
rect 9864 35284 9916 35290
rect 9864 35226 9916 35232
rect 9864 35080 9916 35086
rect 9864 35022 9916 35028
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 9680 33040 9732 33046
rect 9680 32982 9732 32988
rect 9784 32570 9812 33458
rect 9876 33114 9904 35022
rect 10048 34944 10100 34950
rect 10046 34912 10048 34921
rect 10100 34912 10102 34921
rect 10046 34847 10102 34856
rect 10048 34400 10100 34406
rect 10048 34342 10100 34348
rect 10060 34105 10088 34342
rect 10046 34096 10102 34105
rect 10046 34031 10102 34040
rect 10046 33416 10102 33425
rect 10046 33351 10048 33360
rect 10100 33351 10102 33360
rect 10048 33322 10100 33328
rect 9864 33108 9916 33114
rect 9864 33050 9916 33056
rect 10048 32768 10100 32774
rect 10048 32710 10100 32716
rect 10060 32609 10088 32710
rect 10046 32600 10102 32609
rect 9772 32564 9824 32570
rect 10046 32535 10102 32544
rect 9772 32506 9824 32512
rect 9109 32124 9417 32144
rect 9109 32122 9115 32124
rect 9171 32122 9195 32124
rect 9251 32122 9275 32124
rect 9331 32122 9355 32124
rect 9411 32122 9417 32124
rect 9171 32070 9173 32122
rect 9353 32070 9355 32122
rect 9109 32068 9115 32070
rect 9171 32068 9195 32070
rect 9251 32068 9275 32070
rect 9331 32068 9355 32070
rect 9411 32068 9417 32070
rect 9109 32048 9417 32068
rect 10048 31952 10100 31958
rect 10048 31894 10100 31900
rect 10060 31793 10088 31894
rect 10046 31784 10102 31793
rect 10046 31719 10102 31728
rect 10048 31136 10100 31142
rect 10046 31104 10048 31113
rect 10100 31104 10102 31113
rect 9109 31036 9417 31056
rect 10046 31039 10102 31048
rect 9109 31034 9115 31036
rect 9171 31034 9195 31036
rect 9251 31034 9275 31036
rect 9331 31034 9355 31036
rect 9411 31034 9417 31036
rect 9171 30982 9173 31034
rect 9353 30982 9355 31034
rect 9109 30980 9115 30982
rect 9171 30980 9195 30982
rect 9251 30980 9275 30982
rect 9331 30980 9355 30982
rect 9411 30980 9417 30982
rect 9109 30960 9417 30980
rect 9496 30728 9548 30734
rect 9496 30670 9548 30676
rect 9109 29948 9417 29968
rect 9109 29946 9115 29948
rect 9171 29946 9195 29948
rect 9251 29946 9275 29948
rect 9331 29946 9355 29948
rect 9411 29946 9417 29948
rect 9171 29894 9173 29946
rect 9353 29894 9355 29946
rect 9109 29892 9115 29894
rect 9171 29892 9195 29894
rect 9251 29892 9275 29894
rect 9331 29892 9355 29894
rect 9411 29892 9417 29894
rect 9109 29872 9417 29892
rect 9508 29481 9536 30670
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 10060 30297 10088 30534
rect 10046 30288 10102 30297
rect 10046 30223 10102 30232
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 9494 29472 9550 29481
rect 9494 29407 9550 29416
rect 9109 28860 9417 28880
rect 9109 28858 9115 28860
rect 9171 28858 9195 28860
rect 9251 28858 9275 28860
rect 9331 28858 9355 28860
rect 9411 28858 9417 28860
rect 9171 28806 9173 28858
rect 9353 28806 9355 28858
rect 9109 28804 9115 28806
rect 9171 28804 9195 28806
rect 9251 28804 9275 28806
rect 9331 28804 9355 28806
rect 9411 28804 9417 28806
rect 9109 28784 9417 28804
rect 10152 28801 10180 29990
rect 10138 28792 10194 28801
rect 10138 28727 10194 28736
rect 10140 28416 10192 28422
rect 10140 28358 10192 28364
rect 10152 27985 10180 28358
rect 10138 27976 10194 27985
rect 10138 27911 10194 27920
rect 9109 27772 9417 27792
rect 9109 27770 9115 27772
rect 9171 27770 9195 27772
rect 9251 27770 9275 27772
rect 9331 27770 9355 27772
rect 9411 27770 9417 27772
rect 9171 27718 9173 27770
rect 9353 27718 9355 27770
rect 9109 27716 9115 27718
rect 9171 27716 9195 27718
rect 9251 27716 9275 27718
rect 9331 27716 9355 27718
rect 9411 27716 9417 27718
rect 9109 27696 9417 27716
rect 10140 27328 10192 27334
rect 10140 27270 10192 27276
rect 10152 27169 10180 27270
rect 10138 27160 10194 27169
rect 10138 27095 10194 27104
rect 9109 26684 9417 26704
rect 9109 26682 9115 26684
rect 9171 26682 9195 26684
rect 9251 26682 9275 26684
rect 9331 26682 9355 26684
rect 9411 26682 9417 26684
rect 9171 26630 9173 26682
rect 9353 26630 9355 26682
rect 9109 26628 9115 26630
rect 9171 26628 9195 26630
rect 9251 26628 9275 26630
rect 9331 26628 9355 26630
rect 9411 26628 9417 26630
rect 9109 26608 9417 26628
rect 10138 26480 10194 26489
rect 10138 26415 10140 26424
rect 10192 26415 10194 26424
rect 10140 26386 10192 26392
rect 10138 25664 10194 25673
rect 9109 25596 9417 25616
rect 10138 25599 10194 25608
rect 9109 25594 9115 25596
rect 9171 25594 9195 25596
rect 9251 25594 9275 25596
rect 9331 25594 9355 25596
rect 9411 25594 9417 25596
rect 9171 25542 9173 25594
rect 9353 25542 9355 25594
rect 9109 25540 9115 25542
rect 9171 25540 9195 25542
rect 9251 25540 9275 25542
rect 9331 25540 9355 25542
rect 9411 25540 9417 25542
rect 9109 25520 9417 25540
rect 10152 25498 10180 25599
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10138 24848 10194 24857
rect 10138 24783 10140 24792
rect 10192 24783 10194 24792
rect 10140 24754 10192 24760
rect 9109 24508 9417 24528
rect 9109 24506 9115 24508
rect 9171 24506 9195 24508
rect 9251 24506 9275 24508
rect 9331 24506 9355 24508
rect 9411 24506 9417 24508
rect 9171 24454 9173 24506
rect 9353 24454 9355 24506
rect 9109 24452 9115 24454
rect 9171 24452 9195 24454
rect 9251 24452 9275 24454
rect 9331 24452 9355 24454
rect 9411 24452 9417 24454
rect 9109 24432 9417 24452
rect 10138 24168 10194 24177
rect 10138 24103 10194 24112
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9109 23420 9417 23440
rect 9109 23418 9115 23420
rect 9171 23418 9195 23420
rect 9251 23418 9275 23420
rect 9331 23418 9355 23420
rect 9411 23418 9417 23420
rect 9171 23366 9173 23418
rect 9353 23366 9355 23418
rect 9109 23364 9115 23366
rect 9171 23364 9195 23366
rect 9251 23364 9275 23366
rect 9331 23364 9355 23366
rect 9411 23364 9417 23366
rect 9109 23344 9417 23364
rect 9876 23322 9904 23666
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 10060 23361 10088 23462
rect 10046 23352 10102 23361
rect 9864 23316 9916 23322
rect 10152 23322 10180 24103
rect 10046 23287 10102 23296
rect 10140 23316 10192 23322
rect 9864 23258 9916 23264
rect 10140 23258 10192 23264
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9109 22332 9417 22352
rect 9109 22330 9115 22332
rect 9171 22330 9195 22332
rect 9251 22330 9275 22332
rect 9331 22330 9355 22332
rect 9411 22330 9417 22332
rect 9171 22278 9173 22330
rect 9353 22278 9355 22330
rect 9109 22276 9115 22278
rect 9171 22276 9195 22278
rect 9251 22276 9275 22278
rect 9331 22276 9355 22278
rect 9411 22276 9417 22278
rect 9109 22256 9417 22276
rect 9784 21894 9812 22578
rect 10046 22536 10102 22545
rect 10046 22471 10048 22480
rect 10100 22471 10102 22480
rect 10048 22442 10100 22448
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9109 21244 9417 21264
rect 9109 21242 9115 21244
rect 9171 21242 9195 21244
rect 9251 21242 9275 21244
rect 9331 21242 9355 21244
rect 9411 21242 9417 21244
rect 9171 21190 9173 21242
rect 9353 21190 9355 21242
rect 9109 21188 9115 21190
rect 9171 21188 9195 21190
rect 9251 21188 9275 21190
rect 9331 21188 9355 21190
rect 9411 21188 9417 21190
rect 9109 21168 9417 21188
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9109 20156 9417 20176
rect 9109 20154 9115 20156
rect 9171 20154 9195 20156
rect 9251 20154 9275 20156
rect 9331 20154 9355 20156
rect 9411 20154 9417 20156
rect 9171 20102 9173 20154
rect 9353 20102 9355 20154
rect 9109 20100 9115 20102
rect 9171 20100 9195 20102
rect 9251 20100 9275 20102
rect 9331 20100 9355 20102
rect 9411 20100 9417 20102
rect 9109 20080 9417 20100
rect 9109 19068 9417 19088
rect 9109 19066 9115 19068
rect 9171 19066 9195 19068
rect 9251 19066 9275 19068
rect 9331 19066 9355 19068
rect 9411 19066 9417 19068
rect 9171 19014 9173 19066
rect 9353 19014 9355 19066
rect 9109 19012 9115 19014
rect 9171 19012 9195 19014
rect 9251 19012 9275 19014
rect 9331 19012 9355 19014
rect 9411 19012 9417 19014
rect 9109 18992 9417 19012
rect 9692 18426 9720 20402
rect 9784 19514 9812 21490
rect 9876 21146 9904 21966
rect 10048 21888 10100 21894
rect 10046 21856 10048 21865
rect 10100 21856 10102 21865
rect 10046 21791 10102 21800
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 10060 21049 10088 21286
rect 10046 21040 10102 21049
rect 10046 20975 10102 20984
rect 10046 20360 10102 20369
rect 10046 20295 10048 20304
rect 10100 20295 10102 20304
rect 10048 20266 10100 20272
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9876 18970 9904 19790
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 10060 19553 10088 19654
rect 10046 19544 10102 19553
rect 10046 19479 10102 19488
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 10046 18728 10102 18737
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9109 17980 9417 18000
rect 9109 17978 9115 17980
rect 9171 17978 9195 17980
rect 9251 17978 9275 17980
rect 9331 17978 9355 17980
rect 9411 17978 9417 17980
rect 9171 17926 9173 17978
rect 9353 17926 9355 17978
rect 9109 17924 9115 17926
rect 9171 17924 9195 17926
rect 9251 17924 9275 17926
rect 9331 17924 9355 17926
rect 9411 17924 9417 17926
rect 9109 17904 9417 17924
rect 9109 16892 9417 16912
rect 9109 16890 9115 16892
rect 9171 16890 9195 16892
rect 9251 16890 9275 16892
rect 9331 16890 9355 16892
rect 9411 16890 9417 16892
rect 9171 16838 9173 16890
rect 9353 16838 9355 16890
rect 9109 16836 9115 16838
rect 9171 16836 9195 16838
rect 9251 16836 9275 16838
rect 9331 16836 9355 16838
rect 9411 16836 9417 16838
rect 9109 16816 9417 16836
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9109 15804 9417 15824
rect 9109 15802 9115 15804
rect 9171 15802 9195 15804
rect 9251 15802 9275 15804
rect 9331 15802 9355 15804
rect 9411 15802 9417 15804
rect 9171 15750 9173 15802
rect 9353 15750 9355 15802
rect 9109 15748 9115 15750
rect 9171 15748 9195 15750
rect 9251 15748 9275 15750
rect 9331 15748 9355 15750
rect 9411 15748 9417 15750
rect 9109 15728 9417 15748
rect 9109 14716 9417 14736
rect 9109 14714 9115 14716
rect 9171 14714 9195 14716
rect 9251 14714 9275 14716
rect 9331 14714 9355 14716
rect 9411 14714 9417 14716
rect 9171 14662 9173 14714
rect 9353 14662 9355 14714
rect 9109 14660 9115 14662
rect 9171 14660 9195 14662
rect 9251 14660 9275 14662
rect 9331 14660 9355 14662
rect 9411 14660 9417 14662
rect 9109 14640 9417 14660
rect 9692 14074 9720 16526
rect 9784 16454 9812 18702
rect 10046 18663 10102 18672
rect 10060 18630 10088 18663
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9876 15706 9904 17614
rect 9968 17338 9996 18226
rect 10048 18080 10100 18086
rect 10046 18048 10048 18057
rect 10100 18048 10102 18057
rect 10046 17983 10102 17992
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10060 17241 10088 17478
rect 10046 17232 10102 17241
rect 10046 17167 10102 17176
rect 10048 16448 10100 16454
rect 10046 16416 10048 16425
rect 10100 16416 10102 16425
rect 10046 16351 10102 16360
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15745 10088 15846
rect 10046 15736 10102 15745
rect 9864 15700 9916 15706
rect 10046 15671 10102 15680
rect 9864 15642 9916 15648
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10046 14920 10102 14929
rect 10046 14855 10048 14864
rect 10100 14855 10102 14864
rect 10048 14826 10100 14832
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 14113 10088 14214
rect 10046 14104 10102 14113
rect 9680 14068 9732 14074
rect 10046 14039 10102 14048
rect 9680 14010 9732 14016
rect 10152 13870 10180 15438
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 9109 13628 9417 13648
rect 9109 13626 9115 13628
rect 9171 13626 9195 13628
rect 9251 13626 9275 13628
rect 9331 13626 9355 13628
rect 9411 13626 9417 13628
rect 9171 13574 9173 13626
rect 9353 13574 9355 13626
rect 9109 13572 9115 13574
rect 9171 13572 9195 13574
rect 9251 13572 9275 13574
rect 9331 13572 9355 13574
rect 9411 13572 9417 13574
rect 9109 13552 9417 13572
rect 10060 13433 10088 13670
rect 10046 13424 10102 13433
rect 10046 13359 10102 13368
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9109 12540 9417 12560
rect 9109 12538 9115 12540
rect 9171 12538 9195 12540
rect 9251 12538 9275 12540
rect 9331 12538 9355 12540
rect 9411 12538 9417 12540
rect 9171 12486 9173 12538
rect 9353 12486 9355 12538
rect 9109 12484 9115 12486
rect 9171 12484 9195 12486
rect 9251 12484 9275 12486
rect 9331 12484 9355 12486
rect 9411 12484 9417 12486
rect 9109 12464 9417 12484
rect 9784 12102 9812 12786
rect 10048 12640 10100 12646
rect 10046 12608 10048 12617
rect 10100 12608 10102 12617
rect 10046 12543 10102 12552
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9876 11558 9904 12174
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10060 11801 10088 12038
rect 10046 11792 10102 11801
rect 10046 11727 10102 11736
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9109 11452 9417 11472
rect 9109 11450 9115 11452
rect 9171 11450 9195 11452
rect 9251 11450 9275 11452
rect 9331 11450 9355 11452
rect 9411 11450 9417 11452
rect 9171 11398 9173 11450
rect 9353 11398 9355 11450
rect 9109 11396 9115 11398
rect 9171 11396 9195 11398
rect 9251 11396 9275 11398
rect 9331 11396 9355 11398
rect 9411 11396 9417 11398
rect 9109 11376 9417 11396
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9692 10674 9720 11222
rect 10060 11121 10088 11222
rect 10046 11112 10102 11121
rect 9772 11076 9824 11082
rect 10046 11047 10102 11056
rect 9772 11018 9824 11024
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9109 10364 9417 10384
rect 9109 10362 9115 10364
rect 9171 10362 9195 10364
rect 9251 10362 9275 10364
rect 9331 10362 9355 10364
rect 9411 10362 9417 10364
rect 9171 10310 9173 10362
rect 9353 10310 9355 10362
rect 9109 10308 9115 10310
rect 9171 10308 9195 10310
rect 9251 10308 9275 10310
rect 9331 10308 9355 10310
rect 9411 10308 9417 10310
rect 9109 10288 9417 10308
rect 9784 9586 9812 11018
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 10060 10305 10088 10406
rect 10046 10296 10102 10305
rect 10046 10231 10102 10240
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9109 9276 9417 9296
rect 9109 9274 9115 9276
rect 9171 9274 9195 9276
rect 9251 9274 9275 9276
rect 9331 9274 9355 9276
rect 9411 9274 9417 9276
rect 9171 9222 9173 9274
rect 9353 9222 9355 9274
rect 9109 9220 9115 9222
rect 9171 9220 9195 9222
rect 9251 9220 9275 9222
rect 9331 9220 9355 9222
rect 9411 9220 9417 9222
rect 9109 9200 9417 9220
rect 9876 8974 9904 9862
rect 10152 9722 10180 9998
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10046 9480 10102 9489
rect 10046 9415 10048 9424
rect 10100 9415 10102 9424
rect 10048 9386 10100 9392
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 10048 8832 10100 8838
rect 10046 8800 10048 8809
rect 10100 8800 10102 8809
rect 10046 8735 10102 8744
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9109 8188 9417 8208
rect 9109 8186 9115 8188
rect 9171 8186 9195 8188
rect 9251 8186 9275 8188
rect 9331 8186 9355 8188
rect 9411 8186 9417 8188
rect 9171 8134 9173 8186
rect 9353 8134 9355 8186
rect 9109 8132 9115 8134
rect 9171 8132 9195 8134
rect 9251 8132 9275 8134
rect 9331 8132 9355 8134
rect 9411 8132 9417 8134
rect 9109 8112 9417 8132
rect 10060 7993 10088 8230
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9876 7410 9904 7754
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9864 7200 9916 7206
rect 10048 7200 10100 7206
rect 9864 7142 9916 7148
rect 10046 7168 10048 7177
rect 10100 7168 10102 7177
rect 9109 7100 9417 7120
rect 9109 7098 9115 7100
rect 9171 7098 9195 7100
rect 9251 7098 9275 7100
rect 9331 7098 9355 7100
rect 9411 7098 9417 7100
rect 9171 7046 9173 7098
rect 9353 7046 9355 7098
rect 9109 7044 9115 7046
rect 9171 7044 9195 7046
rect 9251 7044 9275 7046
rect 9331 7044 9355 7046
rect 9411 7044 9417 7046
rect 9109 7024 9417 7044
rect 7944 6886 8064 6914
rect 7477 6556 7785 6576
rect 7477 6554 7483 6556
rect 7539 6554 7563 6556
rect 7619 6554 7643 6556
rect 7699 6554 7723 6556
rect 7779 6554 7785 6556
rect 7539 6502 7541 6554
rect 7721 6502 7723 6554
rect 7477 6500 7483 6502
rect 7539 6500 7563 6502
rect 7619 6500 7643 6502
rect 7699 6500 7723 6502
rect 7779 6500 7785 6502
rect 7477 6480 7785 6500
rect 5845 6012 6153 6032
rect 5845 6010 5851 6012
rect 5907 6010 5931 6012
rect 5987 6010 6011 6012
rect 6067 6010 6091 6012
rect 6147 6010 6153 6012
rect 5907 5958 5909 6010
rect 6089 5958 6091 6010
rect 5845 5956 5851 5958
rect 5907 5956 5931 5958
rect 5987 5956 6011 5958
rect 6067 5956 6091 5958
rect 6147 5956 6153 5958
rect 5845 5936 6153 5956
rect 7477 5468 7785 5488
rect 7477 5466 7483 5468
rect 7539 5466 7563 5468
rect 7619 5466 7643 5468
rect 7699 5466 7723 5468
rect 7779 5466 7785 5468
rect 7539 5414 7541 5466
rect 7721 5414 7723 5466
rect 7477 5412 7483 5414
rect 7539 5412 7563 5414
rect 7619 5412 7643 5414
rect 7699 5412 7723 5414
rect 7779 5412 7785 5414
rect 7477 5392 7785 5412
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 5845 4924 6153 4944
rect 5845 4922 5851 4924
rect 5907 4922 5931 4924
rect 5987 4922 6011 4924
rect 6067 4922 6091 4924
rect 6147 4922 6153 4924
rect 5907 4870 5909 4922
rect 6089 4870 6091 4922
rect 5845 4868 5851 4870
rect 5907 4868 5931 4870
rect 5987 4868 6011 4870
rect 6067 4868 6091 4870
rect 6147 4868 6153 4870
rect 5845 4848 6153 4868
rect 7116 4622 7144 4966
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7477 4380 7785 4400
rect 7477 4378 7483 4380
rect 7539 4378 7563 4380
rect 7619 4378 7643 4380
rect 7699 4378 7723 4380
rect 7779 4378 7785 4380
rect 7539 4326 7541 4378
rect 7721 4326 7723 4378
rect 7477 4324 7483 4326
rect 7539 4324 7563 4326
rect 7619 4324 7643 4326
rect 7699 4324 7723 4326
rect 7779 4324 7785 4326
rect 7477 4304 7785 4324
rect 5845 3836 6153 3856
rect 5845 3834 5851 3836
rect 5907 3834 5931 3836
rect 5987 3834 6011 3836
rect 6067 3834 6091 3836
rect 6147 3834 6153 3836
rect 5907 3782 5909 3834
rect 6089 3782 6091 3834
rect 5845 3780 5851 3782
rect 5907 3780 5931 3782
rect 5987 3780 6011 3782
rect 6067 3780 6091 3782
rect 6147 3780 6153 3782
rect 5845 3760 6153 3780
rect 7944 3466 7972 6886
rect 9109 6012 9417 6032
rect 9109 6010 9115 6012
rect 9171 6010 9195 6012
rect 9251 6010 9275 6012
rect 9331 6010 9355 6012
rect 9411 6010 9417 6012
rect 9171 5958 9173 6010
rect 9353 5958 9355 6010
rect 9109 5956 9115 5958
rect 9171 5956 9195 5958
rect 9251 5956 9275 5958
rect 9331 5956 9355 5958
rect 9411 5956 9417 5958
rect 9109 5936 9417 5956
rect 9876 5234 9904 7142
rect 10046 7103 10102 7112
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6497 10088 6598
rect 10046 6488 10102 6497
rect 10046 6423 10102 6432
rect 10046 5672 10102 5681
rect 10046 5607 10102 5616
rect 10060 5574 10088 5607
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9109 4924 9417 4944
rect 9109 4922 9115 4924
rect 9171 4922 9195 4924
rect 9251 4922 9275 4924
rect 9331 4922 9355 4924
rect 9411 4922 9417 4924
rect 9171 4870 9173 4922
rect 9353 4870 9355 4922
rect 9109 4868 9115 4870
rect 9171 4868 9195 4870
rect 9251 4868 9275 4870
rect 9331 4868 9355 4870
rect 9411 4868 9417 4870
rect 9109 4848 9417 4868
rect 10060 4865 10088 4966
rect 10046 4856 10102 4865
rect 9864 4820 9916 4826
rect 10046 4791 10102 4800
rect 9864 4762 9916 4768
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7477 3292 7785 3312
rect 7477 3290 7483 3292
rect 7539 3290 7563 3292
rect 7619 3290 7643 3292
rect 7699 3290 7723 3292
rect 7779 3290 7785 3292
rect 7539 3238 7541 3290
rect 7721 3238 7723 3290
rect 7477 3236 7483 3238
rect 7539 3236 7563 3238
rect 7619 3236 7643 3238
rect 7699 3236 7723 3238
rect 7779 3236 7785 3238
rect 7477 3216 7785 3236
rect 8036 3058 8064 3878
rect 9109 3836 9417 3856
rect 9109 3834 9115 3836
rect 9171 3834 9195 3836
rect 9251 3834 9275 3836
rect 9331 3834 9355 3836
rect 9411 3834 9417 3836
rect 9171 3782 9173 3834
rect 9353 3782 9355 3834
rect 9109 3780 9115 3782
rect 9171 3780 9195 3782
rect 9251 3780 9275 3782
rect 9331 3780 9355 3782
rect 9411 3780 9417 3782
rect 9109 3760 9417 3780
rect 9784 3058 9812 4626
rect 9876 3534 9904 4762
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4185 10088 4422
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10048 3392 10100 3398
rect 10046 3360 10048 3369
rect 10100 3360 10102 3369
rect 10046 3295 10102 3304
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 5845 2748 6153 2768
rect 5845 2746 5851 2748
rect 5907 2746 5931 2748
rect 5987 2746 6011 2748
rect 6067 2746 6091 2748
rect 6147 2746 6153 2748
rect 5907 2694 5909 2746
rect 6089 2694 6091 2746
rect 5845 2692 5851 2694
rect 5907 2692 5931 2694
rect 5987 2692 6011 2694
rect 6067 2692 6091 2694
rect 6147 2692 6153 2694
rect 5845 2672 6153 2692
rect 9109 2748 9417 2768
rect 9109 2746 9115 2748
rect 9171 2746 9195 2748
rect 9251 2746 9275 2748
rect 9331 2746 9355 2748
rect 9411 2746 9417 2748
rect 9171 2694 9173 2746
rect 9353 2694 9355 2746
rect 9109 2692 9115 2694
rect 9171 2692 9195 2694
rect 9251 2692 9275 2694
rect 9331 2692 9355 2694
rect 9411 2692 9417 2694
rect 9109 2672 9417 2692
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 3606 2272 3662 2281
rect 3606 2207 3662 2216
rect 3988 1873 4016 2382
rect 4213 2204 4521 2224
rect 4213 2202 4219 2204
rect 4275 2202 4299 2204
rect 4355 2202 4379 2204
rect 4435 2202 4459 2204
rect 4515 2202 4521 2204
rect 4275 2150 4277 2202
rect 4457 2150 4459 2202
rect 4213 2148 4219 2150
rect 4275 2148 4299 2150
rect 4355 2148 4379 2150
rect 4435 2148 4459 2150
rect 4515 2148 4521 2150
rect 4213 2128 4521 2148
rect 3974 1864 4030 1873
rect 3974 1799 4030 1808
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 2872 1080 2924 1086
rect 2870 1048 2872 1057
rect 2924 1048 2926 1057
rect 2870 983 2926 992
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 2780 536 2832 542
rect 2780 478 2832 484
rect 2792 241 2820 478
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 2962 0 3018 800
rect 4632 542 4660 2382
rect 5276 1086 5304 2382
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 7477 2204 7785 2224
rect 7477 2202 7483 2204
rect 7539 2202 7563 2204
rect 7619 2202 7643 2204
rect 7699 2202 7723 2204
rect 7779 2202 7785 2204
rect 7539 2150 7541 2202
rect 7721 2150 7723 2202
rect 7477 2148 7483 2150
rect 7539 2148 7563 2150
rect 7619 2148 7643 2150
rect 7699 2148 7723 2150
rect 7779 2148 7785 2150
rect 7477 2128 7785 2148
rect 5264 1080 5316 1086
rect 5264 1022 5316 1028
rect 4620 536 4672 542
rect 4620 478 4672 484
rect 8942 0 8998 800
rect 9324 377 9352 2246
rect 9508 1873 9536 2790
rect 9876 2446 9904 2858
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2553 10088 2790
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 9494 1864 9550 1873
rect 9494 1799 9550 1808
rect 10060 1057 10088 2246
rect 10046 1048 10102 1057
rect 10046 983 10102 992
rect 9310 368 9366 377
rect 9310 303 9366 312
<< via2 >>
rect 2962 79600 3018 79656
rect 1398 79192 1454 79248
rect 2778 78784 2834 78840
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 10046 79464 10102 79520
rect 3514 78376 3570 78432
rect 3422 77560 3478 77616
rect 1490 74432 1546 74488
rect 1398 74296 1454 74352
rect 1398 73208 1454 73264
rect 1398 71848 1454 71904
rect 1214 71032 1270 71088
rect 1306 70624 1362 70680
rect 1398 70216 1454 70272
rect 1306 68720 1362 68776
rect 1398 68040 1454 68096
rect 1306 67632 1362 67688
rect 1398 67224 1454 67280
rect 1398 66816 1454 66872
rect 1398 66272 1454 66328
rect 1398 65864 1454 65920
rect 2042 72392 2098 72448
rect 1766 66408 1822 66464
rect 1674 66156 1730 66192
rect 1674 66136 1676 66156
rect 1676 66136 1728 66156
rect 1728 66136 1730 66156
rect 1766 65628 1768 65648
rect 1768 65628 1820 65648
rect 1820 65628 1822 65648
rect 1398 62464 1454 62520
rect 1766 65592 1822 65628
rect 1490 62056 1546 62112
rect 1490 61684 1492 61704
rect 1492 61684 1544 61704
rect 1544 61684 1546 61704
rect 1490 61648 1546 61684
rect 1398 61104 1454 61160
rect 1490 60696 1546 60752
rect 1398 59880 1454 59936
rect 1398 59064 1454 59120
rect 1582 58792 1638 58848
rect 1490 58520 1546 58576
rect 1490 56888 1546 56944
rect 1490 56480 1546 56536
rect 1490 55392 1546 55448
rect 1674 58540 1730 58576
rect 1674 58520 1676 58540
rect 1676 58520 1728 58540
rect 1728 58520 1730 58540
rect 1398 55256 1454 55312
rect 1398 53896 1454 53952
rect 1490 53488 1546 53544
rect 1398 52128 1454 52184
rect 2226 71440 2282 71496
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 2962 76200 3018 76256
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 2778 73616 2834 73672
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2134 64912 2190 64968
rect 2226 63724 2228 63744
rect 2228 63724 2280 63744
rect 2280 63724 2282 63744
rect 2226 63688 2282 63724
rect 2778 72800 2834 72856
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 3330 76472 3386 76528
rect 4066 77968 4122 78024
rect 3146 75792 3202 75848
rect 3146 74976 3202 75032
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 2962 69808 3018 69864
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 2870 68756 2872 68776
rect 2872 68756 2924 68776
rect 2924 68756 2926 68776
rect 2870 68720 2926 68756
rect 3054 68856 3110 68912
rect 2962 68448 3018 68504
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 3330 69264 3386 69320
rect 3606 75384 3662 75440
rect 4219 77274 4275 77276
rect 4299 77274 4355 77276
rect 4379 77274 4435 77276
rect 4459 77274 4515 77276
rect 4219 77222 4265 77274
rect 4265 77222 4275 77274
rect 4299 77222 4329 77274
rect 4329 77222 4341 77274
rect 4341 77222 4355 77274
rect 4379 77222 4393 77274
rect 4393 77222 4405 77274
rect 4405 77222 4435 77274
rect 4459 77222 4469 77274
rect 4469 77222 4515 77274
rect 4219 77220 4275 77222
rect 4299 77220 4355 77222
rect 4379 77220 4435 77222
rect 4459 77220 4515 77222
rect 3974 77016 4030 77072
rect 9494 77968 9550 78024
rect 5851 77818 5907 77820
rect 5931 77818 5987 77820
rect 6011 77818 6067 77820
rect 6091 77818 6147 77820
rect 5851 77766 5897 77818
rect 5897 77766 5907 77818
rect 5931 77766 5961 77818
rect 5961 77766 5973 77818
rect 5973 77766 5987 77818
rect 6011 77766 6025 77818
rect 6025 77766 6037 77818
rect 6037 77766 6067 77818
rect 6091 77766 6101 77818
rect 6101 77766 6147 77818
rect 5851 77764 5907 77766
rect 5931 77764 5987 77766
rect 6011 77764 6067 77766
rect 6091 77764 6147 77766
rect 9115 77818 9171 77820
rect 9195 77818 9251 77820
rect 9275 77818 9331 77820
rect 9355 77818 9411 77820
rect 9115 77766 9161 77818
rect 9161 77766 9171 77818
rect 9195 77766 9225 77818
rect 9225 77766 9237 77818
rect 9237 77766 9251 77818
rect 9275 77766 9289 77818
rect 9289 77766 9301 77818
rect 9301 77766 9331 77818
rect 9355 77766 9365 77818
rect 9365 77766 9411 77818
rect 9115 77764 9171 77766
rect 9195 77764 9251 77766
rect 9275 77764 9331 77766
rect 9355 77764 9411 77766
rect 7483 77274 7539 77276
rect 7563 77274 7619 77276
rect 7643 77274 7699 77276
rect 7723 77274 7779 77276
rect 7483 77222 7529 77274
rect 7529 77222 7539 77274
rect 7563 77222 7593 77274
rect 7593 77222 7605 77274
rect 7605 77222 7619 77274
rect 7643 77222 7657 77274
rect 7657 77222 7669 77274
rect 7669 77222 7699 77274
rect 7723 77222 7733 77274
rect 7733 77222 7779 77274
rect 7483 77220 7539 77222
rect 7563 77220 7619 77222
rect 7643 77220 7699 77222
rect 7723 77220 7779 77222
rect 9402 77152 9458 77208
rect 10966 78668 11022 78704
rect 10966 78648 10968 78668
rect 10968 78648 11020 78668
rect 11020 78648 11022 78668
rect 4219 76186 4275 76188
rect 4299 76186 4355 76188
rect 4379 76186 4435 76188
rect 4459 76186 4515 76188
rect 4219 76134 4265 76186
rect 4265 76134 4275 76186
rect 4299 76134 4329 76186
rect 4329 76134 4341 76186
rect 4341 76134 4355 76186
rect 4379 76134 4393 76186
rect 4393 76134 4405 76186
rect 4405 76134 4435 76186
rect 4459 76134 4469 76186
rect 4469 76134 4515 76186
rect 4219 76132 4275 76134
rect 4299 76132 4355 76134
rect 4379 76132 4435 76134
rect 4459 76132 4515 76134
rect 2962 65456 3018 65512
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 2778 64268 2780 64288
rect 2780 64268 2832 64288
rect 2832 64268 2834 64288
rect 2778 64232 2834 64268
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 3054 63280 3110 63336
rect 2870 62872 2926 62928
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 2502 60832 2558 60888
rect 2502 60696 2558 60752
rect 2318 58520 2374 58576
rect 2778 60580 2834 60616
rect 2778 60560 2780 60580
rect 2780 60560 2832 60580
rect 2832 60560 2834 60580
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2502 60152 2558 60208
rect 2410 58112 2466 58168
rect 2226 57316 2282 57352
rect 2226 57296 2228 57316
rect 2228 57296 2280 57316
rect 2280 57296 2282 57316
rect 2226 55936 2282 55992
rect 1674 51856 1730 51912
rect 1490 51720 1546 51776
rect 1398 50360 1454 50416
rect 1490 49952 1546 50008
rect 1214 40160 1270 40216
rect 1214 38800 1270 38856
rect 1490 48320 1546 48376
rect 1490 47776 1546 47832
rect 1490 47540 1492 47560
rect 1492 47540 1544 47560
rect 1544 47540 1546 47560
rect 1490 47504 1546 47540
rect 1490 46960 1546 47016
rect 1490 46552 1546 46608
rect 1490 46144 1546 46200
rect 1582 45872 1638 45928
rect 1490 45772 1492 45792
rect 1492 45772 1544 45792
rect 1544 45772 1546 45792
rect 1490 45736 1546 45772
rect 1490 44784 1546 44840
rect 1490 41384 1546 41440
rect 1490 39616 1546 39672
rect 1490 37712 1546 37768
rect 1490 37032 1546 37088
rect 1490 35808 1546 35864
rect 1490 34992 1546 35048
rect 1950 48320 2006 48376
rect 1858 45056 1914 45112
rect 2318 55564 2320 55584
rect 2320 55564 2372 55584
rect 2372 55564 2374 55584
rect 2318 55528 2374 55564
rect 2318 52536 2374 52592
rect 2226 50904 2282 50960
rect 2686 59628 2742 59664
rect 2686 59608 2688 59628
rect 2688 59608 2740 59628
rect 2740 59608 2742 59628
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2778 57740 2780 57760
rect 2780 57740 2832 57760
rect 2832 57740 2834 57760
rect 2778 57704 2834 57740
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 3054 59492 3110 59528
rect 3054 59472 3056 59492
rect 3056 59472 3108 59492
rect 3108 59472 3110 59492
rect 3054 57876 3056 57896
rect 3056 57876 3108 57896
rect 3108 57876 3110 57896
rect 3054 57840 3110 57876
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 2778 54304 2834 54360
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 3054 52964 3110 53000
rect 3054 52944 3056 52964
rect 3056 52944 3108 52964
rect 3108 52944 3110 52964
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 3054 51312 3110 51368
rect 2410 49580 2412 49600
rect 2412 49580 2464 49600
rect 2464 49580 2466 49600
rect 2410 49544 2466 49580
rect 2226 49136 2282 49192
rect 2226 45328 2282 45384
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2778 48728 2834 48784
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2962 48272 3018 48328
rect 2778 47776 2834 47832
rect 2686 47504 2742 47560
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 2778 46416 2834 46472
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 2778 44956 2780 44976
rect 2780 44956 2832 44976
rect 2832 44956 2834 44976
rect 2318 43560 2374 43616
rect 2778 44920 2834 44956
rect 2778 44376 2834 44432
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 2962 43832 3018 43888
rect 3330 65048 3386 65104
rect 2778 43152 2834 43208
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2226 41792 2282 41848
rect 1950 40840 2006 40896
rect 1490 32408 1546 32464
rect 1582 31864 1638 31920
rect 1490 31048 1546 31104
rect 1490 30640 1546 30696
rect 2226 40568 2282 40624
rect 2134 40024 2190 40080
rect 2962 42608 3018 42664
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2226 37032 2282 37088
rect 2226 36760 2282 36816
rect 1858 31864 1914 31920
rect 1858 31728 1914 31784
rect 1214 22072 1270 22128
rect 1398 28056 1454 28112
rect 1398 26288 1454 26344
rect 1490 25064 1546 25120
rect 1398 24248 1454 24304
rect 1490 22888 1546 22944
rect 1398 21120 1454 21176
rect 1766 28056 1822 28112
rect 2318 36216 2374 36272
rect 2594 41112 2650 41168
rect 3054 42200 3110 42256
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 3054 40996 3110 41032
rect 3054 40976 3056 40996
rect 3056 40976 3108 40996
rect 3108 40976 3110 40996
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 2778 39244 2780 39264
rect 2780 39244 2832 39264
rect 2832 39244 2834 39264
rect 2778 39208 2834 39244
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 2962 37984 3018 38040
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 3054 36644 3110 36680
rect 3054 36624 3056 36644
rect 3056 36624 3108 36644
rect 3108 36624 3110 36644
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 3054 35556 3110 35592
rect 3054 35536 3056 35556
rect 3056 35536 3108 35556
rect 3108 35536 3110 35556
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 2410 34040 2466 34096
rect 2318 33632 2374 33688
rect 2318 33260 2320 33280
rect 2320 33260 2372 33280
rect 2372 33260 2374 33280
rect 2318 33224 2374 33260
rect 2318 32816 2374 32872
rect 2042 27512 2098 27568
rect 1490 16496 1546 16552
rect 1398 15544 1454 15600
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 3514 56888 3570 56944
rect 3514 47796 3570 47832
rect 3514 47776 3516 47796
rect 3516 47776 3568 47796
rect 3568 47776 3570 47796
rect 3882 64504 3938 64560
rect 3698 50360 3754 50416
rect 3698 47096 3754 47152
rect 3422 45328 3478 45384
rect 3422 41520 3478 41576
rect 3330 41112 3386 41168
rect 3238 37304 3294 37360
rect 3238 34448 3294 34504
rect 4219 75098 4275 75100
rect 4299 75098 4355 75100
rect 4379 75098 4435 75100
rect 4459 75098 4515 75100
rect 4219 75046 4265 75098
rect 4265 75046 4275 75098
rect 4299 75046 4329 75098
rect 4329 75046 4341 75098
rect 4341 75046 4355 75098
rect 4379 75046 4393 75098
rect 4393 75046 4405 75098
rect 4405 75046 4435 75098
rect 4459 75046 4469 75098
rect 4469 75046 4515 75098
rect 4219 75044 4275 75046
rect 4299 75044 4355 75046
rect 4379 75044 4435 75046
rect 4459 75044 4515 75046
rect 4219 74010 4275 74012
rect 4299 74010 4355 74012
rect 4379 74010 4435 74012
rect 4459 74010 4515 74012
rect 4219 73958 4265 74010
rect 4265 73958 4275 74010
rect 4299 73958 4329 74010
rect 4329 73958 4341 74010
rect 4341 73958 4355 74010
rect 4379 73958 4393 74010
rect 4393 73958 4405 74010
rect 4405 73958 4435 74010
rect 4459 73958 4469 74010
rect 4469 73958 4515 74010
rect 4219 73956 4275 73958
rect 4299 73956 4355 73958
rect 4379 73956 4435 73958
rect 4459 73956 4515 73958
rect 4219 72922 4275 72924
rect 4299 72922 4355 72924
rect 4379 72922 4435 72924
rect 4459 72922 4515 72924
rect 4219 72870 4265 72922
rect 4265 72870 4275 72922
rect 4299 72870 4329 72922
rect 4329 72870 4341 72922
rect 4341 72870 4355 72922
rect 4379 72870 4393 72922
rect 4393 72870 4405 72922
rect 4405 72870 4435 72922
rect 4459 72870 4469 72922
rect 4469 72870 4515 72922
rect 4219 72868 4275 72870
rect 4299 72868 4355 72870
rect 4379 72868 4435 72870
rect 4459 72868 4515 72870
rect 4219 71834 4275 71836
rect 4299 71834 4355 71836
rect 4379 71834 4435 71836
rect 4459 71834 4515 71836
rect 4219 71782 4265 71834
rect 4265 71782 4275 71834
rect 4299 71782 4329 71834
rect 4329 71782 4341 71834
rect 4341 71782 4355 71834
rect 4379 71782 4393 71834
rect 4393 71782 4405 71834
rect 4405 71782 4435 71834
rect 4459 71782 4469 71834
rect 4469 71782 4515 71834
rect 4219 71780 4275 71782
rect 4299 71780 4355 71782
rect 4379 71780 4435 71782
rect 4459 71780 4515 71782
rect 4219 70746 4275 70748
rect 4299 70746 4355 70748
rect 4379 70746 4435 70748
rect 4459 70746 4515 70748
rect 4219 70694 4265 70746
rect 4265 70694 4275 70746
rect 4299 70694 4329 70746
rect 4329 70694 4341 70746
rect 4341 70694 4355 70746
rect 4379 70694 4393 70746
rect 4393 70694 4405 70746
rect 4405 70694 4435 70746
rect 4459 70694 4469 70746
rect 4469 70694 4515 70746
rect 4219 70692 4275 70694
rect 4299 70692 4355 70694
rect 4379 70692 4435 70694
rect 4459 70692 4515 70694
rect 4219 69658 4275 69660
rect 4299 69658 4355 69660
rect 4379 69658 4435 69660
rect 4459 69658 4515 69660
rect 4219 69606 4265 69658
rect 4265 69606 4275 69658
rect 4299 69606 4329 69658
rect 4329 69606 4341 69658
rect 4341 69606 4355 69658
rect 4379 69606 4393 69658
rect 4393 69606 4405 69658
rect 4405 69606 4435 69658
rect 4459 69606 4469 69658
rect 4469 69606 4515 69658
rect 4219 69604 4275 69606
rect 4299 69604 4355 69606
rect 4379 69604 4435 69606
rect 4459 69604 4515 69606
rect 4219 68570 4275 68572
rect 4299 68570 4355 68572
rect 4379 68570 4435 68572
rect 4459 68570 4515 68572
rect 4219 68518 4265 68570
rect 4265 68518 4275 68570
rect 4299 68518 4329 68570
rect 4329 68518 4341 68570
rect 4341 68518 4355 68570
rect 4379 68518 4393 68570
rect 4393 68518 4405 68570
rect 4405 68518 4435 68570
rect 4459 68518 4469 68570
rect 4469 68518 4515 68570
rect 4219 68516 4275 68518
rect 4299 68516 4355 68518
rect 4379 68516 4435 68518
rect 4459 68516 4515 68518
rect 4219 67482 4275 67484
rect 4299 67482 4355 67484
rect 4379 67482 4435 67484
rect 4459 67482 4515 67484
rect 4219 67430 4265 67482
rect 4265 67430 4275 67482
rect 4299 67430 4329 67482
rect 4329 67430 4341 67482
rect 4341 67430 4355 67482
rect 4379 67430 4393 67482
rect 4393 67430 4405 67482
rect 4405 67430 4435 67482
rect 4459 67430 4469 67482
rect 4469 67430 4515 67482
rect 4219 67428 4275 67430
rect 4299 67428 4355 67430
rect 4379 67428 4435 67430
rect 4459 67428 4515 67430
rect 4219 66394 4275 66396
rect 4299 66394 4355 66396
rect 4379 66394 4435 66396
rect 4459 66394 4515 66396
rect 4219 66342 4265 66394
rect 4265 66342 4275 66394
rect 4299 66342 4329 66394
rect 4329 66342 4341 66394
rect 4341 66342 4355 66394
rect 4379 66342 4393 66394
rect 4393 66342 4405 66394
rect 4405 66342 4435 66394
rect 4459 66342 4469 66394
rect 4469 66342 4515 66394
rect 4219 66340 4275 66342
rect 4299 66340 4355 66342
rect 4379 66340 4435 66342
rect 4459 66340 4515 66342
rect 4219 65306 4275 65308
rect 4299 65306 4355 65308
rect 4379 65306 4435 65308
rect 4459 65306 4515 65308
rect 4219 65254 4265 65306
rect 4265 65254 4275 65306
rect 4299 65254 4329 65306
rect 4329 65254 4341 65306
rect 4341 65254 4355 65306
rect 4379 65254 4393 65306
rect 4393 65254 4405 65306
rect 4405 65254 4435 65306
rect 4459 65254 4469 65306
rect 4469 65254 4515 65306
rect 4219 65252 4275 65254
rect 4299 65252 4355 65254
rect 4379 65252 4435 65254
rect 4459 65252 4515 65254
rect 4219 64218 4275 64220
rect 4299 64218 4355 64220
rect 4379 64218 4435 64220
rect 4459 64218 4515 64220
rect 4219 64166 4265 64218
rect 4265 64166 4275 64218
rect 4299 64166 4329 64218
rect 4329 64166 4341 64218
rect 4341 64166 4355 64218
rect 4379 64166 4393 64218
rect 4393 64166 4405 64218
rect 4405 64166 4435 64218
rect 4459 64166 4469 64218
rect 4469 64166 4515 64218
rect 4219 64164 4275 64166
rect 4299 64164 4355 64166
rect 4379 64164 4435 64166
rect 4459 64164 4515 64166
rect 4219 63130 4275 63132
rect 4299 63130 4355 63132
rect 4379 63130 4435 63132
rect 4459 63130 4515 63132
rect 4219 63078 4265 63130
rect 4265 63078 4275 63130
rect 4299 63078 4329 63130
rect 4329 63078 4341 63130
rect 4341 63078 4355 63130
rect 4379 63078 4393 63130
rect 4393 63078 4405 63130
rect 4405 63078 4435 63130
rect 4459 63078 4469 63130
rect 4469 63078 4515 63130
rect 4219 63076 4275 63078
rect 4299 63076 4355 63078
rect 4379 63076 4435 63078
rect 4459 63076 4515 63078
rect 4219 62042 4275 62044
rect 4299 62042 4355 62044
rect 4379 62042 4435 62044
rect 4459 62042 4515 62044
rect 4219 61990 4265 62042
rect 4265 61990 4275 62042
rect 4299 61990 4329 62042
rect 4329 61990 4341 62042
rect 4341 61990 4355 62042
rect 4379 61990 4393 62042
rect 4393 61990 4405 62042
rect 4405 61990 4435 62042
rect 4459 61990 4469 62042
rect 4469 61990 4515 62042
rect 4219 61988 4275 61990
rect 4299 61988 4355 61990
rect 4379 61988 4435 61990
rect 4459 61988 4515 61990
rect 4219 60954 4275 60956
rect 4299 60954 4355 60956
rect 4379 60954 4435 60956
rect 4459 60954 4515 60956
rect 4219 60902 4265 60954
rect 4265 60902 4275 60954
rect 4299 60902 4329 60954
rect 4329 60902 4341 60954
rect 4341 60902 4355 60954
rect 4379 60902 4393 60954
rect 4393 60902 4405 60954
rect 4405 60902 4435 60954
rect 4459 60902 4469 60954
rect 4469 60902 4515 60954
rect 4219 60900 4275 60902
rect 4299 60900 4355 60902
rect 4379 60900 4435 60902
rect 4459 60900 4515 60902
rect 4219 59866 4275 59868
rect 4299 59866 4355 59868
rect 4379 59866 4435 59868
rect 4459 59866 4515 59868
rect 4219 59814 4265 59866
rect 4265 59814 4275 59866
rect 4299 59814 4329 59866
rect 4329 59814 4341 59866
rect 4341 59814 4355 59866
rect 4379 59814 4393 59866
rect 4393 59814 4405 59866
rect 4405 59814 4435 59866
rect 4459 59814 4469 59866
rect 4469 59814 4515 59866
rect 4219 59812 4275 59814
rect 4299 59812 4355 59814
rect 4379 59812 4435 59814
rect 4459 59812 4515 59814
rect 4219 58778 4275 58780
rect 4299 58778 4355 58780
rect 4379 58778 4435 58780
rect 4459 58778 4515 58780
rect 4219 58726 4265 58778
rect 4265 58726 4275 58778
rect 4299 58726 4329 58778
rect 4329 58726 4341 58778
rect 4341 58726 4355 58778
rect 4379 58726 4393 58778
rect 4393 58726 4405 58778
rect 4405 58726 4435 58778
rect 4459 58726 4469 58778
rect 4469 58726 4515 58778
rect 4219 58724 4275 58726
rect 4299 58724 4355 58726
rect 4379 58724 4435 58726
rect 4459 58724 4515 58726
rect 4219 57690 4275 57692
rect 4299 57690 4355 57692
rect 4379 57690 4435 57692
rect 4459 57690 4515 57692
rect 4219 57638 4265 57690
rect 4265 57638 4275 57690
rect 4299 57638 4329 57690
rect 4329 57638 4341 57690
rect 4341 57638 4355 57690
rect 4379 57638 4393 57690
rect 4393 57638 4405 57690
rect 4405 57638 4435 57690
rect 4459 57638 4469 57690
rect 4469 57638 4515 57690
rect 4219 57636 4275 57638
rect 4299 57636 4355 57638
rect 4379 57636 4435 57638
rect 4459 57636 4515 57638
rect 4219 56602 4275 56604
rect 4299 56602 4355 56604
rect 4379 56602 4435 56604
rect 4459 56602 4515 56604
rect 4219 56550 4265 56602
rect 4265 56550 4275 56602
rect 4299 56550 4329 56602
rect 4329 56550 4341 56602
rect 4341 56550 4355 56602
rect 4379 56550 4393 56602
rect 4393 56550 4405 56602
rect 4405 56550 4435 56602
rect 4459 56550 4469 56602
rect 4469 56550 4515 56602
rect 4219 56548 4275 56550
rect 4299 56548 4355 56550
rect 4379 56548 4435 56550
rect 4459 56548 4515 56550
rect 4219 55514 4275 55516
rect 4299 55514 4355 55516
rect 4379 55514 4435 55516
rect 4459 55514 4515 55516
rect 4219 55462 4265 55514
rect 4265 55462 4275 55514
rect 4299 55462 4329 55514
rect 4329 55462 4341 55514
rect 4341 55462 4355 55514
rect 4379 55462 4393 55514
rect 4393 55462 4405 55514
rect 4405 55462 4435 55514
rect 4459 55462 4469 55514
rect 4469 55462 4515 55514
rect 4219 55460 4275 55462
rect 4299 55460 4355 55462
rect 4379 55460 4435 55462
rect 4459 55460 4515 55462
rect 4219 54426 4275 54428
rect 4299 54426 4355 54428
rect 4379 54426 4435 54428
rect 4459 54426 4515 54428
rect 4219 54374 4265 54426
rect 4265 54374 4275 54426
rect 4299 54374 4329 54426
rect 4329 54374 4341 54426
rect 4341 54374 4355 54426
rect 4379 54374 4393 54426
rect 4393 54374 4405 54426
rect 4405 54374 4435 54426
rect 4459 54374 4469 54426
rect 4469 54374 4515 54426
rect 4219 54372 4275 54374
rect 4299 54372 4355 54374
rect 4379 54372 4435 54374
rect 4459 54372 4515 54374
rect 4219 53338 4275 53340
rect 4299 53338 4355 53340
rect 4379 53338 4435 53340
rect 4459 53338 4515 53340
rect 4219 53286 4265 53338
rect 4265 53286 4275 53338
rect 4299 53286 4329 53338
rect 4329 53286 4341 53338
rect 4341 53286 4355 53338
rect 4379 53286 4393 53338
rect 4393 53286 4405 53338
rect 4405 53286 4435 53338
rect 4459 53286 4469 53338
rect 4469 53286 4515 53338
rect 4219 53284 4275 53286
rect 4299 53284 4355 53286
rect 4379 53284 4435 53286
rect 4459 53284 4515 53286
rect 4219 52250 4275 52252
rect 4299 52250 4355 52252
rect 4379 52250 4435 52252
rect 4459 52250 4515 52252
rect 4219 52198 4265 52250
rect 4265 52198 4275 52250
rect 4299 52198 4329 52250
rect 4329 52198 4341 52250
rect 4341 52198 4355 52250
rect 4379 52198 4393 52250
rect 4393 52198 4405 52250
rect 4405 52198 4435 52250
rect 4459 52198 4469 52250
rect 4469 52198 4515 52250
rect 4219 52196 4275 52198
rect 4299 52196 4355 52198
rect 4379 52196 4435 52198
rect 4459 52196 4515 52198
rect 4219 51162 4275 51164
rect 4299 51162 4355 51164
rect 4379 51162 4435 51164
rect 4459 51162 4515 51164
rect 4219 51110 4265 51162
rect 4265 51110 4275 51162
rect 4299 51110 4329 51162
rect 4329 51110 4341 51162
rect 4341 51110 4355 51162
rect 4379 51110 4393 51162
rect 4393 51110 4405 51162
rect 4405 51110 4435 51162
rect 4459 51110 4469 51162
rect 4469 51110 4515 51162
rect 4219 51108 4275 51110
rect 4299 51108 4355 51110
rect 4379 51108 4435 51110
rect 4459 51108 4515 51110
rect 4618 50360 4674 50416
rect 4219 50074 4275 50076
rect 4299 50074 4355 50076
rect 4379 50074 4435 50076
rect 4459 50074 4515 50076
rect 4219 50022 4265 50074
rect 4265 50022 4275 50074
rect 4299 50022 4329 50074
rect 4329 50022 4341 50074
rect 4341 50022 4355 50074
rect 4379 50022 4393 50074
rect 4393 50022 4405 50074
rect 4405 50022 4435 50074
rect 4459 50022 4469 50074
rect 4469 50022 4515 50074
rect 4219 50020 4275 50022
rect 4299 50020 4355 50022
rect 4379 50020 4435 50022
rect 4459 50020 4515 50022
rect 3606 41384 3662 41440
rect 3422 38392 3478 38448
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 2778 31456 2834 31512
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 3606 38292 3608 38312
rect 3608 38292 3660 38312
rect 3660 38292 3662 38312
rect 3606 38256 3662 38292
rect 3514 33496 3570 33552
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 3146 28736 3202 28792
rect 3238 28600 3294 28656
rect 2870 28500 2872 28520
rect 2872 28500 2924 28520
rect 2924 28500 2926 28520
rect 2870 28464 2926 28500
rect 2410 27648 2466 27704
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 2962 27240 3018 27296
rect 3146 26832 3202 26888
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 3054 25880 3110 25936
rect 2870 25744 2926 25800
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2778 24656 2834 24712
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 2962 23160 3018 23216
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 3146 21664 3202 21720
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 2778 20304 2834 20360
rect 1674 13504 1730 13560
rect 1398 12280 1454 12336
rect 1306 11736 1362 11792
rect 1398 11328 1454 11384
rect 1858 12552 1914 12608
rect 1306 10920 1362 10976
rect 1398 10376 1454 10432
rect 1306 9968 1362 10024
rect 1398 9560 1454 9616
rect 1398 9152 1454 9208
rect 1398 7384 1454 7440
rect 1398 6568 1454 6624
rect 1398 4800 1454 4856
rect 1306 3576 1362 3632
rect 1398 3168 1454 3224
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2962 19896 3018 19952
rect 2778 19216 2834 19272
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 3146 19488 3202 19544
rect 2962 18128 3018 18184
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 2870 17040 2926 17096
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 2226 14728 2282 14784
rect 2778 15952 2834 16008
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 2870 15136 2926 15192
rect 2042 6976 2098 7032
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 3146 13912 3202 13968
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 2778 12960 2834 13016
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 2042 5208 2098 5264
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 4219 48986 4275 48988
rect 4299 48986 4355 48988
rect 4379 48986 4435 48988
rect 4459 48986 4515 48988
rect 4219 48934 4265 48986
rect 4265 48934 4275 48986
rect 4299 48934 4329 48986
rect 4329 48934 4341 48986
rect 4341 48934 4355 48986
rect 4379 48934 4393 48986
rect 4393 48934 4405 48986
rect 4405 48934 4435 48986
rect 4459 48934 4469 48986
rect 4469 48934 4515 48986
rect 4219 48932 4275 48934
rect 4299 48932 4355 48934
rect 4379 48932 4435 48934
rect 4459 48932 4515 48934
rect 4526 48728 4582 48784
rect 4219 47898 4275 47900
rect 4299 47898 4355 47900
rect 4379 47898 4435 47900
rect 4459 47898 4515 47900
rect 4219 47846 4265 47898
rect 4265 47846 4275 47898
rect 4299 47846 4329 47898
rect 4329 47846 4341 47898
rect 4341 47846 4355 47898
rect 4379 47846 4393 47898
rect 4393 47846 4405 47898
rect 4405 47846 4435 47898
rect 4459 47846 4469 47898
rect 4469 47846 4515 47898
rect 4219 47844 4275 47846
rect 4299 47844 4355 47846
rect 4379 47844 4435 47846
rect 4459 47844 4515 47846
rect 4219 46810 4275 46812
rect 4299 46810 4355 46812
rect 4379 46810 4435 46812
rect 4459 46810 4515 46812
rect 4219 46758 4265 46810
rect 4265 46758 4275 46810
rect 4299 46758 4329 46810
rect 4329 46758 4341 46810
rect 4341 46758 4355 46810
rect 4379 46758 4393 46810
rect 4393 46758 4405 46810
rect 4405 46758 4435 46810
rect 4459 46758 4469 46810
rect 4469 46758 4515 46810
rect 4219 46756 4275 46758
rect 4299 46756 4355 46758
rect 4379 46756 4435 46758
rect 4459 46756 4515 46758
rect 4434 46008 4490 46064
rect 4219 45722 4275 45724
rect 4299 45722 4355 45724
rect 4379 45722 4435 45724
rect 4459 45722 4515 45724
rect 4219 45670 4265 45722
rect 4265 45670 4275 45722
rect 4299 45670 4329 45722
rect 4329 45670 4341 45722
rect 4341 45670 4355 45722
rect 4379 45670 4393 45722
rect 4393 45670 4405 45722
rect 4405 45670 4435 45722
rect 4459 45670 4469 45722
rect 4469 45670 4515 45722
rect 4219 45668 4275 45670
rect 4299 45668 4355 45670
rect 4379 45668 4435 45670
rect 4459 45668 4515 45670
rect 3974 41384 4030 41440
rect 4219 44634 4275 44636
rect 4299 44634 4355 44636
rect 4379 44634 4435 44636
rect 4459 44634 4515 44636
rect 4219 44582 4265 44634
rect 4265 44582 4275 44634
rect 4299 44582 4329 44634
rect 4329 44582 4341 44634
rect 4341 44582 4355 44634
rect 4379 44582 4393 44634
rect 4393 44582 4405 44634
rect 4405 44582 4435 44634
rect 4459 44582 4469 44634
rect 4469 44582 4515 44634
rect 4219 44580 4275 44582
rect 4299 44580 4355 44582
rect 4379 44580 4435 44582
rect 4459 44580 4515 44582
rect 4158 44396 4214 44432
rect 4158 44376 4160 44396
rect 4160 44376 4212 44396
rect 4212 44376 4214 44396
rect 4219 43546 4275 43548
rect 4299 43546 4355 43548
rect 4379 43546 4435 43548
rect 4459 43546 4515 43548
rect 4219 43494 4265 43546
rect 4265 43494 4275 43546
rect 4299 43494 4329 43546
rect 4329 43494 4341 43546
rect 4341 43494 4355 43546
rect 4379 43494 4393 43546
rect 4393 43494 4405 43546
rect 4405 43494 4435 43546
rect 4459 43494 4469 43546
rect 4469 43494 4515 43546
rect 4219 43492 4275 43494
rect 4299 43492 4355 43494
rect 4379 43492 4435 43494
rect 4459 43492 4515 43494
rect 4219 42458 4275 42460
rect 4299 42458 4355 42460
rect 4379 42458 4435 42460
rect 4459 42458 4515 42460
rect 4219 42406 4265 42458
rect 4265 42406 4275 42458
rect 4299 42406 4329 42458
rect 4329 42406 4341 42458
rect 4341 42406 4355 42458
rect 4379 42406 4393 42458
rect 4393 42406 4405 42458
rect 4405 42406 4435 42458
rect 4459 42406 4469 42458
rect 4469 42406 4515 42458
rect 4219 42404 4275 42406
rect 4299 42404 4355 42406
rect 4379 42404 4435 42406
rect 4459 42404 4515 42406
rect 4219 41370 4275 41372
rect 4299 41370 4355 41372
rect 4379 41370 4435 41372
rect 4459 41370 4515 41372
rect 4219 41318 4265 41370
rect 4265 41318 4275 41370
rect 4299 41318 4329 41370
rect 4329 41318 4341 41370
rect 4341 41318 4355 41370
rect 4379 41318 4393 41370
rect 4393 41318 4405 41370
rect 4405 41318 4435 41370
rect 4459 41318 4469 41370
rect 4469 41318 4515 41370
rect 4219 41316 4275 41318
rect 4299 41316 4355 41318
rect 4379 41316 4435 41318
rect 4459 41316 4515 41318
rect 4219 40282 4275 40284
rect 4299 40282 4355 40284
rect 4379 40282 4435 40284
rect 4459 40282 4515 40284
rect 4219 40230 4265 40282
rect 4265 40230 4275 40282
rect 4299 40230 4329 40282
rect 4329 40230 4341 40282
rect 4341 40230 4355 40282
rect 4379 40230 4393 40282
rect 4393 40230 4405 40282
rect 4405 40230 4435 40282
rect 4459 40230 4469 40282
rect 4469 40230 4515 40282
rect 4219 40228 4275 40230
rect 4299 40228 4355 40230
rect 4379 40228 4435 40230
rect 4459 40228 4515 40230
rect 4219 39194 4275 39196
rect 4299 39194 4355 39196
rect 4379 39194 4435 39196
rect 4459 39194 4515 39196
rect 4219 39142 4265 39194
rect 4265 39142 4275 39194
rect 4299 39142 4329 39194
rect 4329 39142 4341 39194
rect 4341 39142 4355 39194
rect 4379 39142 4393 39194
rect 4393 39142 4405 39194
rect 4405 39142 4435 39194
rect 4459 39142 4469 39194
rect 4469 39142 4515 39194
rect 4219 39140 4275 39142
rect 4299 39140 4355 39142
rect 4379 39140 4435 39142
rect 4459 39140 4515 39142
rect 4219 38106 4275 38108
rect 4299 38106 4355 38108
rect 4379 38106 4435 38108
rect 4459 38106 4515 38108
rect 4219 38054 4265 38106
rect 4265 38054 4275 38106
rect 4299 38054 4329 38106
rect 4329 38054 4341 38106
rect 4341 38054 4355 38106
rect 4379 38054 4393 38106
rect 4393 38054 4405 38106
rect 4405 38054 4435 38106
rect 4459 38054 4469 38106
rect 4469 38054 4515 38106
rect 4219 38052 4275 38054
rect 4299 38052 4355 38054
rect 4379 38052 4435 38054
rect 4459 38052 4515 38054
rect 4219 37018 4275 37020
rect 4299 37018 4355 37020
rect 4379 37018 4435 37020
rect 4459 37018 4515 37020
rect 4219 36966 4265 37018
rect 4265 36966 4275 37018
rect 4299 36966 4329 37018
rect 4329 36966 4341 37018
rect 4341 36966 4355 37018
rect 4379 36966 4393 37018
rect 4393 36966 4405 37018
rect 4405 36966 4435 37018
rect 4459 36966 4469 37018
rect 4469 36966 4515 37018
rect 4219 36964 4275 36966
rect 4299 36964 4355 36966
rect 4379 36964 4435 36966
rect 4459 36964 4515 36966
rect 4219 35930 4275 35932
rect 4299 35930 4355 35932
rect 4379 35930 4435 35932
rect 4459 35930 4515 35932
rect 4219 35878 4265 35930
rect 4265 35878 4275 35930
rect 4299 35878 4329 35930
rect 4329 35878 4341 35930
rect 4341 35878 4355 35930
rect 4379 35878 4393 35930
rect 4393 35878 4405 35930
rect 4405 35878 4435 35930
rect 4459 35878 4469 35930
rect 4469 35878 4515 35930
rect 4219 35876 4275 35878
rect 4299 35876 4355 35878
rect 4379 35876 4435 35878
rect 4459 35876 4515 35878
rect 5170 45464 5226 45520
rect 5078 42472 5134 42528
rect 4219 34842 4275 34844
rect 4299 34842 4355 34844
rect 4379 34842 4435 34844
rect 4459 34842 4515 34844
rect 4219 34790 4265 34842
rect 4265 34790 4275 34842
rect 4299 34790 4329 34842
rect 4329 34790 4341 34842
rect 4341 34790 4355 34842
rect 4379 34790 4393 34842
rect 4393 34790 4405 34842
rect 4405 34790 4435 34842
rect 4459 34790 4469 34842
rect 4469 34790 4515 34842
rect 4219 34788 4275 34790
rect 4299 34788 4355 34790
rect 4379 34788 4435 34790
rect 4459 34788 4515 34790
rect 4219 33754 4275 33756
rect 4299 33754 4355 33756
rect 4379 33754 4435 33756
rect 4459 33754 4515 33756
rect 4219 33702 4265 33754
rect 4265 33702 4275 33754
rect 4299 33702 4329 33754
rect 4329 33702 4341 33754
rect 4341 33702 4355 33754
rect 4379 33702 4393 33754
rect 4393 33702 4405 33754
rect 4405 33702 4435 33754
rect 4459 33702 4469 33754
rect 4469 33702 4515 33754
rect 4219 33700 4275 33702
rect 4299 33700 4355 33702
rect 4379 33700 4435 33702
rect 4459 33700 4515 33702
rect 3790 32000 3846 32056
rect 3974 30232 4030 30288
rect 3790 30096 3846 30152
rect 3422 22480 3478 22536
rect 3882 29688 3938 29744
rect 3974 29280 4030 29336
rect 3974 23704 4030 23760
rect 3422 17720 3478 17776
rect 3054 8744 3110 8800
rect 3606 21936 3662 21992
rect 4219 32666 4275 32668
rect 4299 32666 4355 32668
rect 4379 32666 4435 32668
rect 4459 32666 4515 32668
rect 4219 32614 4265 32666
rect 4265 32614 4275 32666
rect 4299 32614 4329 32666
rect 4329 32614 4341 32666
rect 4341 32614 4355 32666
rect 4379 32614 4393 32666
rect 4393 32614 4405 32666
rect 4405 32614 4435 32666
rect 4459 32614 4469 32666
rect 4469 32614 4515 32666
rect 4219 32612 4275 32614
rect 4299 32612 4355 32614
rect 4379 32612 4435 32614
rect 4459 32612 4515 32614
rect 4219 31578 4275 31580
rect 4299 31578 4355 31580
rect 4379 31578 4435 31580
rect 4459 31578 4515 31580
rect 4219 31526 4265 31578
rect 4265 31526 4275 31578
rect 4299 31526 4329 31578
rect 4329 31526 4341 31578
rect 4341 31526 4355 31578
rect 4379 31526 4393 31578
rect 4393 31526 4405 31578
rect 4405 31526 4435 31578
rect 4459 31526 4469 31578
rect 4469 31526 4515 31578
rect 4219 31524 4275 31526
rect 4299 31524 4355 31526
rect 4379 31524 4435 31526
rect 4459 31524 4515 31526
rect 4219 30490 4275 30492
rect 4299 30490 4355 30492
rect 4379 30490 4435 30492
rect 4459 30490 4515 30492
rect 4219 30438 4265 30490
rect 4265 30438 4275 30490
rect 4299 30438 4329 30490
rect 4329 30438 4341 30490
rect 4341 30438 4355 30490
rect 4379 30438 4393 30490
rect 4393 30438 4405 30490
rect 4405 30438 4435 30490
rect 4459 30438 4469 30490
rect 4469 30438 4515 30490
rect 4219 30436 4275 30438
rect 4299 30436 4355 30438
rect 4379 30436 4435 30438
rect 4459 30436 4515 30438
rect 4219 29402 4275 29404
rect 4299 29402 4355 29404
rect 4379 29402 4435 29404
rect 4459 29402 4515 29404
rect 4219 29350 4265 29402
rect 4265 29350 4275 29402
rect 4299 29350 4329 29402
rect 4329 29350 4341 29402
rect 4341 29350 4355 29402
rect 4379 29350 4393 29402
rect 4393 29350 4405 29402
rect 4405 29350 4435 29402
rect 4459 29350 4469 29402
rect 4469 29350 4515 29402
rect 4219 29348 4275 29350
rect 4299 29348 4355 29350
rect 4379 29348 4435 29350
rect 4459 29348 4515 29350
rect 4219 28314 4275 28316
rect 4299 28314 4355 28316
rect 4379 28314 4435 28316
rect 4459 28314 4515 28316
rect 4219 28262 4265 28314
rect 4265 28262 4275 28314
rect 4299 28262 4329 28314
rect 4329 28262 4341 28314
rect 4341 28262 4355 28314
rect 4379 28262 4393 28314
rect 4393 28262 4405 28314
rect 4405 28262 4435 28314
rect 4459 28262 4469 28314
rect 4469 28262 4515 28314
rect 4219 28260 4275 28262
rect 4299 28260 4355 28262
rect 4379 28260 4435 28262
rect 4459 28260 4515 28262
rect 4219 27226 4275 27228
rect 4299 27226 4355 27228
rect 4379 27226 4435 27228
rect 4459 27226 4515 27228
rect 4219 27174 4265 27226
rect 4265 27174 4275 27226
rect 4299 27174 4329 27226
rect 4329 27174 4341 27226
rect 4341 27174 4355 27226
rect 4379 27174 4393 27226
rect 4393 27174 4405 27226
rect 4405 27174 4435 27226
rect 4459 27174 4469 27226
rect 4469 27174 4515 27226
rect 4219 27172 4275 27174
rect 4299 27172 4355 27174
rect 4379 27172 4435 27174
rect 4459 27172 4515 27174
rect 4219 26138 4275 26140
rect 4299 26138 4355 26140
rect 4379 26138 4435 26140
rect 4459 26138 4515 26140
rect 4219 26086 4265 26138
rect 4265 26086 4275 26138
rect 4299 26086 4329 26138
rect 4329 26086 4341 26138
rect 4341 26086 4355 26138
rect 4379 26086 4393 26138
rect 4393 26086 4405 26138
rect 4405 26086 4435 26138
rect 4459 26086 4469 26138
rect 4469 26086 4515 26138
rect 4219 26084 4275 26086
rect 4299 26084 4355 26086
rect 4379 26084 4435 26086
rect 4459 26084 4515 26086
rect 4219 25050 4275 25052
rect 4299 25050 4355 25052
rect 4379 25050 4435 25052
rect 4459 25050 4515 25052
rect 4219 24998 4265 25050
rect 4265 24998 4275 25050
rect 4299 24998 4329 25050
rect 4329 24998 4341 25050
rect 4341 24998 4355 25050
rect 4379 24998 4393 25050
rect 4393 24998 4405 25050
rect 4405 24998 4435 25050
rect 4459 24998 4469 25050
rect 4469 24998 4515 25050
rect 4219 24996 4275 24998
rect 4299 24996 4355 24998
rect 4379 24996 4435 24998
rect 4459 24996 4515 24998
rect 4219 23962 4275 23964
rect 4299 23962 4355 23964
rect 4379 23962 4435 23964
rect 4459 23962 4515 23964
rect 4219 23910 4265 23962
rect 4265 23910 4275 23962
rect 4299 23910 4329 23962
rect 4329 23910 4341 23962
rect 4341 23910 4355 23962
rect 4379 23910 4393 23962
rect 4393 23910 4405 23962
rect 4405 23910 4435 23962
rect 4459 23910 4469 23962
rect 4469 23910 4515 23962
rect 4219 23908 4275 23910
rect 4299 23908 4355 23910
rect 4379 23908 4435 23910
rect 4459 23908 4515 23910
rect 4219 22874 4275 22876
rect 4299 22874 4355 22876
rect 4379 22874 4435 22876
rect 4459 22874 4515 22876
rect 4219 22822 4265 22874
rect 4265 22822 4275 22874
rect 4299 22822 4329 22874
rect 4329 22822 4341 22874
rect 4341 22822 4355 22874
rect 4379 22822 4393 22874
rect 4393 22822 4405 22874
rect 4405 22822 4435 22874
rect 4459 22822 4469 22874
rect 4469 22822 4515 22874
rect 4219 22820 4275 22822
rect 4299 22820 4355 22822
rect 4379 22820 4435 22822
rect 4459 22820 4515 22822
rect 4219 21786 4275 21788
rect 4299 21786 4355 21788
rect 4379 21786 4435 21788
rect 4459 21786 4515 21788
rect 4219 21734 4265 21786
rect 4265 21734 4275 21786
rect 4299 21734 4329 21786
rect 4329 21734 4341 21786
rect 4341 21734 4355 21786
rect 4379 21734 4393 21786
rect 4393 21734 4405 21786
rect 4405 21734 4435 21786
rect 4459 21734 4469 21786
rect 4469 21734 4515 21786
rect 4219 21732 4275 21734
rect 4299 21732 4355 21734
rect 4379 21732 4435 21734
rect 4459 21732 4515 21734
rect 3974 20712 4030 20768
rect 4219 20698 4275 20700
rect 4299 20698 4355 20700
rect 4379 20698 4435 20700
rect 4459 20698 4515 20700
rect 4219 20646 4265 20698
rect 4265 20646 4275 20698
rect 4299 20646 4329 20698
rect 4329 20646 4341 20698
rect 4341 20646 4355 20698
rect 4379 20646 4393 20698
rect 4393 20646 4405 20698
rect 4405 20646 4435 20698
rect 4459 20646 4469 20698
rect 4469 20646 4515 20698
rect 4219 20644 4275 20646
rect 4299 20644 4355 20646
rect 4379 20644 4435 20646
rect 4459 20644 4515 20646
rect 4219 19610 4275 19612
rect 4299 19610 4355 19612
rect 4379 19610 4435 19612
rect 4459 19610 4515 19612
rect 4219 19558 4265 19610
rect 4265 19558 4275 19610
rect 4299 19558 4329 19610
rect 4329 19558 4341 19610
rect 4341 19558 4355 19610
rect 4379 19558 4393 19610
rect 4393 19558 4405 19610
rect 4405 19558 4435 19610
rect 4459 19558 4469 19610
rect 4469 19558 4515 19610
rect 4219 19556 4275 19558
rect 4299 19556 4355 19558
rect 4379 19556 4435 19558
rect 4459 19556 4515 19558
rect 3974 18536 4030 18592
rect 3974 17312 4030 17368
rect 3974 14356 3976 14376
rect 3976 14356 4028 14376
rect 4028 14356 4030 14376
rect 3974 14320 4030 14356
rect 3514 8336 3570 8392
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 2962 5752 3018 5808
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 3330 6160 3386 6216
rect 4219 18522 4275 18524
rect 4299 18522 4355 18524
rect 4379 18522 4435 18524
rect 4459 18522 4515 18524
rect 4219 18470 4265 18522
rect 4265 18470 4275 18522
rect 4299 18470 4329 18522
rect 4329 18470 4341 18522
rect 4341 18470 4355 18522
rect 4379 18470 4393 18522
rect 4393 18470 4405 18522
rect 4405 18470 4435 18522
rect 4459 18470 4469 18522
rect 4469 18470 4515 18522
rect 4219 18468 4275 18470
rect 4299 18468 4355 18470
rect 4379 18468 4435 18470
rect 4459 18468 4515 18470
rect 4219 17434 4275 17436
rect 4299 17434 4355 17436
rect 4379 17434 4435 17436
rect 4459 17434 4515 17436
rect 4219 17382 4265 17434
rect 4265 17382 4275 17434
rect 4299 17382 4329 17434
rect 4329 17382 4341 17434
rect 4341 17382 4355 17434
rect 4379 17382 4393 17434
rect 4393 17382 4405 17434
rect 4405 17382 4435 17434
rect 4459 17382 4469 17434
rect 4469 17382 4515 17434
rect 4219 17380 4275 17382
rect 4299 17380 4355 17382
rect 4379 17380 4435 17382
rect 4459 17380 4515 17382
rect 4219 16346 4275 16348
rect 4299 16346 4355 16348
rect 4379 16346 4435 16348
rect 4459 16346 4515 16348
rect 4219 16294 4265 16346
rect 4265 16294 4275 16346
rect 4299 16294 4329 16346
rect 4329 16294 4341 16346
rect 4341 16294 4355 16346
rect 4379 16294 4393 16346
rect 4393 16294 4405 16346
rect 4405 16294 4435 16346
rect 4459 16294 4469 16346
rect 4469 16294 4515 16346
rect 4219 16292 4275 16294
rect 4299 16292 4355 16294
rect 4379 16292 4435 16294
rect 4459 16292 4515 16294
rect 4219 15258 4275 15260
rect 4299 15258 4355 15260
rect 4379 15258 4435 15260
rect 4459 15258 4515 15260
rect 4219 15206 4265 15258
rect 4265 15206 4275 15258
rect 4299 15206 4329 15258
rect 4329 15206 4341 15258
rect 4341 15206 4355 15258
rect 4379 15206 4393 15258
rect 4393 15206 4405 15258
rect 4405 15206 4435 15258
rect 4459 15206 4469 15258
rect 4469 15206 4515 15258
rect 4219 15204 4275 15206
rect 4299 15204 4355 15206
rect 4379 15204 4435 15206
rect 4459 15204 4515 15206
rect 4219 14170 4275 14172
rect 4299 14170 4355 14172
rect 4379 14170 4435 14172
rect 4459 14170 4515 14172
rect 4219 14118 4265 14170
rect 4265 14118 4275 14170
rect 4299 14118 4329 14170
rect 4329 14118 4341 14170
rect 4341 14118 4355 14170
rect 4379 14118 4393 14170
rect 4393 14118 4405 14170
rect 4405 14118 4435 14170
rect 4459 14118 4469 14170
rect 4469 14118 4515 14170
rect 4219 14116 4275 14118
rect 4299 14116 4355 14118
rect 4379 14116 4435 14118
rect 4459 14116 4515 14118
rect 4219 13082 4275 13084
rect 4299 13082 4355 13084
rect 4379 13082 4435 13084
rect 4459 13082 4515 13084
rect 4219 13030 4265 13082
rect 4265 13030 4275 13082
rect 4299 13030 4329 13082
rect 4329 13030 4341 13082
rect 4341 13030 4355 13082
rect 4379 13030 4393 13082
rect 4393 13030 4405 13082
rect 4405 13030 4435 13082
rect 4459 13030 4469 13082
rect 4469 13030 4515 13082
rect 4219 13028 4275 13030
rect 4299 13028 4355 13030
rect 4379 13028 4435 13030
rect 4459 13028 4515 13030
rect 4219 11994 4275 11996
rect 4299 11994 4355 11996
rect 4379 11994 4435 11996
rect 4459 11994 4515 11996
rect 4219 11942 4265 11994
rect 4265 11942 4275 11994
rect 4299 11942 4329 11994
rect 4329 11942 4341 11994
rect 4341 11942 4355 11994
rect 4379 11942 4393 11994
rect 4393 11942 4405 11994
rect 4405 11942 4435 11994
rect 4459 11942 4469 11994
rect 4469 11942 4515 11994
rect 4219 11940 4275 11942
rect 4299 11940 4355 11942
rect 4379 11940 4435 11942
rect 4459 11940 4515 11942
rect 3790 7828 3792 7848
rect 3792 7828 3844 7848
rect 3844 7828 3846 7848
rect 3790 7792 3846 7828
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 4219 10906 4275 10908
rect 4299 10906 4355 10908
rect 4379 10906 4435 10908
rect 4459 10906 4515 10908
rect 4219 10854 4265 10906
rect 4265 10854 4275 10906
rect 4299 10854 4329 10906
rect 4329 10854 4341 10906
rect 4341 10854 4355 10906
rect 4379 10854 4393 10906
rect 4393 10854 4405 10906
rect 4405 10854 4435 10906
rect 4459 10854 4469 10906
rect 4469 10854 4515 10906
rect 4219 10852 4275 10854
rect 4299 10852 4355 10854
rect 4379 10852 4435 10854
rect 4459 10852 4515 10854
rect 4219 9818 4275 9820
rect 4299 9818 4355 9820
rect 4379 9818 4435 9820
rect 4459 9818 4515 9820
rect 4219 9766 4265 9818
rect 4265 9766 4275 9818
rect 4299 9766 4329 9818
rect 4329 9766 4341 9818
rect 4341 9766 4355 9818
rect 4379 9766 4393 9818
rect 4393 9766 4405 9818
rect 4405 9766 4435 9818
rect 4459 9766 4469 9818
rect 4469 9766 4515 9818
rect 4219 9764 4275 9766
rect 4299 9764 4355 9766
rect 4379 9764 4435 9766
rect 4459 9764 4515 9766
rect 4219 8730 4275 8732
rect 4299 8730 4355 8732
rect 4379 8730 4435 8732
rect 4459 8730 4515 8732
rect 4219 8678 4265 8730
rect 4265 8678 4275 8730
rect 4299 8678 4329 8730
rect 4329 8678 4341 8730
rect 4341 8678 4355 8730
rect 4379 8678 4393 8730
rect 4393 8678 4405 8730
rect 4405 8678 4435 8730
rect 4459 8678 4469 8730
rect 4469 8678 4515 8730
rect 4219 8676 4275 8678
rect 4299 8676 4355 8678
rect 4379 8676 4435 8678
rect 4459 8676 4515 8678
rect 4219 7642 4275 7644
rect 4299 7642 4355 7644
rect 4379 7642 4435 7644
rect 4459 7642 4515 7644
rect 4219 7590 4265 7642
rect 4265 7590 4275 7642
rect 4299 7590 4329 7642
rect 4329 7590 4341 7642
rect 4341 7590 4355 7642
rect 4379 7590 4393 7642
rect 4393 7590 4405 7642
rect 4405 7590 4435 7642
rect 4459 7590 4469 7642
rect 4469 7590 4515 7642
rect 4219 7588 4275 7590
rect 4299 7588 4355 7590
rect 4379 7588 4435 7590
rect 4459 7588 4515 7590
rect 4219 6554 4275 6556
rect 4299 6554 4355 6556
rect 4379 6554 4435 6556
rect 4459 6554 4515 6556
rect 4219 6502 4265 6554
rect 4265 6502 4275 6554
rect 4299 6502 4329 6554
rect 4329 6502 4341 6554
rect 4341 6502 4355 6554
rect 4379 6502 4393 6554
rect 4393 6502 4405 6554
rect 4405 6502 4435 6554
rect 4459 6502 4469 6554
rect 4469 6502 4515 6554
rect 4219 6500 4275 6502
rect 4299 6500 4355 6502
rect 4379 6500 4435 6502
rect 4459 6500 4515 6502
rect 4219 5466 4275 5468
rect 4299 5466 4355 5468
rect 4379 5466 4435 5468
rect 4459 5466 4515 5468
rect 4219 5414 4265 5466
rect 4265 5414 4275 5466
rect 4299 5414 4329 5466
rect 4329 5414 4341 5466
rect 4341 5414 4355 5466
rect 4379 5414 4393 5466
rect 4393 5414 4405 5466
rect 4405 5414 4435 5466
rect 4459 5414 4469 5466
rect 4469 5414 4515 5466
rect 4219 5412 4275 5414
rect 4299 5412 4355 5414
rect 4379 5412 4435 5414
rect 4459 5412 4515 5414
rect 5851 76730 5907 76732
rect 5931 76730 5987 76732
rect 6011 76730 6067 76732
rect 6091 76730 6147 76732
rect 5851 76678 5897 76730
rect 5897 76678 5907 76730
rect 5931 76678 5961 76730
rect 5961 76678 5973 76730
rect 5973 76678 5987 76730
rect 6011 76678 6025 76730
rect 6025 76678 6037 76730
rect 6037 76678 6067 76730
rect 6091 76678 6101 76730
rect 6101 76678 6147 76730
rect 5851 76676 5907 76678
rect 5931 76676 5987 76678
rect 6011 76676 6067 76678
rect 6091 76676 6147 76678
rect 9115 76730 9171 76732
rect 9195 76730 9251 76732
rect 9275 76730 9331 76732
rect 9355 76730 9411 76732
rect 9115 76678 9161 76730
rect 9161 76678 9171 76730
rect 9195 76678 9225 76730
rect 9225 76678 9237 76730
rect 9237 76678 9251 76730
rect 9275 76678 9289 76730
rect 9289 76678 9301 76730
rect 9301 76678 9331 76730
rect 9355 76678 9365 76730
rect 9365 76678 9411 76730
rect 9115 76676 9171 76678
rect 9195 76676 9251 76678
rect 9275 76676 9331 76678
rect 9355 76676 9411 76678
rect 10138 76372 10140 76392
rect 10140 76372 10192 76392
rect 10192 76372 10194 76392
rect 10138 76336 10194 76372
rect 7483 76186 7539 76188
rect 7563 76186 7619 76188
rect 7643 76186 7699 76188
rect 7723 76186 7779 76188
rect 7483 76134 7529 76186
rect 7529 76134 7539 76186
rect 7563 76134 7593 76186
rect 7593 76134 7605 76186
rect 7605 76134 7619 76186
rect 7643 76134 7657 76186
rect 7657 76134 7669 76186
rect 7669 76134 7699 76186
rect 7723 76134 7733 76186
rect 7733 76134 7779 76186
rect 7483 76132 7539 76134
rect 7563 76132 7619 76134
rect 7643 76132 7699 76134
rect 7723 76132 7779 76134
rect 5851 75642 5907 75644
rect 5931 75642 5987 75644
rect 6011 75642 6067 75644
rect 6091 75642 6147 75644
rect 5851 75590 5897 75642
rect 5897 75590 5907 75642
rect 5931 75590 5961 75642
rect 5961 75590 5973 75642
rect 5973 75590 5987 75642
rect 6011 75590 6025 75642
rect 6025 75590 6037 75642
rect 6037 75590 6067 75642
rect 6091 75590 6101 75642
rect 6101 75590 6147 75642
rect 5851 75588 5907 75590
rect 5931 75588 5987 75590
rect 6011 75588 6067 75590
rect 6091 75588 6147 75590
rect 9115 75642 9171 75644
rect 9195 75642 9251 75644
rect 9275 75642 9331 75644
rect 9355 75642 9411 75644
rect 9115 75590 9161 75642
rect 9161 75590 9171 75642
rect 9195 75590 9225 75642
rect 9225 75590 9237 75642
rect 9237 75590 9251 75642
rect 9275 75590 9289 75642
rect 9289 75590 9301 75642
rect 9301 75590 9331 75642
rect 9355 75590 9365 75642
rect 9365 75590 9411 75642
rect 9115 75588 9171 75590
rect 9195 75588 9251 75590
rect 9275 75588 9331 75590
rect 9355 75588 9411 75590
rect 7483 75098 7539 75100
rect 7563 75098 7619 75100
rect 7643 75098 7699 75100
rect 7723 75098 7779 75100
rect 7483 75046 7529 75098
rect 7529 75046 7539 75098
rect 7563 75046 7593 75098
rect 7593 75046 7605 75098
rect 7605 75046 7619 75098
rect 7643 75046 7657 75098
rect 7657 75046 7669 75098
rect 7669 75046 7699 75098
rect 7723 75046 7733 75098
rect 7733 75046 7779 75098
rect 7483 75044 7539 75046
rect 7563 75044 7619 75046
rect 7643 75044 7699 75046
rect 7723 75044 7779 75046
rect 5851 74554 5907 74556
rect 5931 74554 5987 74556
rect 6011 74554 6067 74556
rect 6091 74554 6147 74556
rect 5851 74502 5897 74554
rect 5897 74502 5907 74554
rect 5931 74502 5961 74554
rect 5961 74502 5973 74554
rect 5973 74502 5987 74554
rect 6011 74502 6025 74554
rect 6025 74502 6037 74554
rect 6037 74502 6067 74554
rect 6091 74502 6101 74554
rect 6101 74502 6147 74554
rect 5851 74500 5907 74502
rect 5931 74500 5987 74502
rect 6011 74500 6067 74502
rect 6091 74500 6147 74502
rect 7483 74010 7539 74012
rect 7563 74010 7619 74012
rect 7643 74010 7699 74012
rect 7723 74010 7779 74012
rect 7483 73958 7529 74010
rect 7529 73958 7539 74010
rect 7563 73958 7593 74010
rect 7593 73958 7605 74010
rect 7605 73958 7619 74010
rect 7643 73958 7657 74010
rect 7657 73958 7669 74010
rect 7669 73958 7699 74010
rect 7723 73958 7733 74010
rect 7733 73958 7779 74010
rect 7483 73956 7539 73958
rect 7563 73956 7619 73958
rect 7643 73956 7699 73958
rect 7723 73956 7779 73958
rect 5851 73466 5907 73468
rect 5931 73466 5987 73468
rect 6011 73466 6067 73468
rect 6091 73466 6147 73468
rect 5851 73414 5897 73466
rect 5897 73414 5907 73466
rect 5931 73414 5961 73466
rect 5961 73414 5973 73466
rect 5973 73414 5987 73466
rect 6011 73414 6025 73466
rect 6025 73414 6037 73466
rect 6037 73414 6067 73466
rect 6091 73414 6101 73466
rect 6101 73414 6147 73466
rect 5851 73412 5907 73414
rect 5931 73412 5987 73414
rect 6011 73412 6067 73414
rect 6091 73412 6147 73414
rect 7483 72922 7539 72924
rect 7563 72922 7619 72924
rect 7643 72922 7699 72924
rect 7723 72922 7779 72924
rect 7483 72870 7529 72922
rect 7529 72870 7539 72922
rect 7563 72870 7593 72922
rect 7593 72870 7605 72922
rect 7605 72870 7619 72922
rect 7643 72870 7657 72922
rect 7657 72870 7669 72922
rect 7669 72870 7699 72922
rect 7723 72870 7733 72922
rect 7733 72870 7779 72922
rect 7483 72868 7539 72870
rect 7563 72868 7619 72870
rect 7643 72868 7699 72870
rect 7723 72868 7779 72870
rect 5851 72378 5907 72380
rect 5931 72378 5987 72380
rect 6011 72378 6067 72380
rect 6091 72378 6147 72380
rect 5851 72326 5897 72378
rect 5897 72326 5907 72378
rect 5931 72326 5961 72378
rect 5961 72326 5973 72378
rect 5973 72326 5987 72378
rect 6011 72326 6025 72378
rect 6025 72326 6037 72378
rect 6037 72326 6067 72378
rect 6091 72326 6101 72378
rect 6101 72326 6147 72378
rect 5851 72324 5907 72326
rect 5931 72324 5987 72326
rect 6011 72324 6067 72326
rect 6091 72324 6147 72326
rect 7483 71834 7539 71836
rect 7563 71834 7619 71836
rect 7643 71834 7699 71836
rect 7723 71834 7779 71836
rect 7483 71782 7529 71834
rect 7529 71782 7539 71834
rect 7563 71782 7593 71834
rect 7593 71782 7605 71834
rect 7605 71782 7619 71834
rect 7643 71782 7657 71834
rect 7657 71782 7669 71834
rect 7669 71782 7699 71834
rect 7723 71782 7733 71834
rect 7733 71782 7779 71834
rect 7483 71780 7539 71782
rect 7563 71780 7619 71782
rect 7643 71780 7699 71782
rect 7723 71780 7779 71782
rect 5851 71290 5907 71292
rect 5931 71290 5987 71292
rect 6011 71290 6067 71292
rect 6091 71290 6147 71292
rect 5851 71238 5897 71290
rect 5897 71238 5907 71290
rect 5931 71238 5961 71290
rect 5961 71238 5973 71290
rect 5973 71238 5987 71290
rect 6011 71238 6025 71290
rect 6025 71238 6037 71290
rect 6037 71238 6067 71290
rect 6091 71238 6101 71290
rect 6101 71238 6147 71290
rect 5851 71236 5907 71238
rect 5931 71236 5987 71238
rect 6011 71236 6067 71238
rect 6091 71236 6147 71238
rect 7483 70746 7539 70748
rect 7563 70746 7619 70748
rect 7643 70746 7699 70748
rect 7723 70746 7779 70748
rect 7483 70694 7529 70746
rect 7529 70694 7539 70746
rect 7563 70694 7593 70746
rect 7593 70694 7605 70746
rect 7605 70694 7619 70746
rect 7643 70694 7657 70746
rect 7657 70694 7669 70746
rect 7669 70694 7699 70746
rect 7723 70694 7733 70746
rect 7733 70694 7779 70746
rect 7483 70692 7539 70694
rect 7563 70692 7619 70694
rect 7643 70692 7699 70694
rect 7723 70692 7779 70694
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 3974 4392 4030 4448
rect 4219 4378 4275 4380
rect 4299 4378 4355 4380
rect 4379 4378 4435 4380
rect 4459 4378 4515 4380
rect 4219 4326 4265 4378
rect 4265 4326 4275 4378
rect 4299 4326 4329 4378
rect 4329 4326 4341 4378
rect 4341 4326 4355 4378
rect 4379 4326 4393 4378
rect 4393 4326 4405 4378
rect 4405 4326 4435 4378
rect 4459 4326 4469 4378
rect 4469 4326 4515 4378
rect 4219 4324 4275 4326
rect 4299 4324 4355 4326
rect 4379 4324 4435 4326
rect 4459 4324 4515 4326
rect 3974 3984 4030 4040
rect 4219 3290 4275 3292
rect 4299 3290 4355 3292
rect 4379 3290 4435 3292
rect 4459 3290 4515 3292
rect 4219 3238 4265 3290
rect 4265 3238 4275 3290
rect 4299 3238 4329 3290
rect 4329 3238 4341 3290
rect 4341 3238 4355 3290
rect 4379 3238 4393 3290
rect 4393 3238 4405 3290
rect 4405 3238 4435 3290
rect 4459 3238 4469 3290
rect 4469 3238 4515 3290
rect 4219 3236 4275 3238
rect 4299 3236 4355 3238
rect 4379 3236 4435 3238
rect 4459 3236 4515 3238
rect 4066 2488 4122 2544
rect 5851 70202 5907 70204
rect 5931 70202 5987 70204
rect 6011 70202 6067 70204
rect 6091 70202 6147 70204
rect 5851 70150 5897 70202
rect 5897 70150 5907 70202
rect 5931 70150 5961 70202
rect 5961 70150 5973 70202
rect 5973 70150 5987 70202
rect 6011 70150 6025 70202
rect 6025 70150 6037 70202
rect 6037 70150 6067 70202
rect 6091 70150 6101 70202
rect 6101 70150 6147 70202
rect 5851 70148 5907 70150
rect 5931 70148 5987 70150
rect 6011 70148 6067 70150
rect 6091 70148 6147 70150
rect 7483 69658 7539 69660
rect 7563 69658 7619 69660
rect 7643 69658 7699 69660
rect 7723 69658 7779 69660
rect 7483 69606 7529 69658
rect 7529 69606 7539 69658
rect 7563 69606 7593 69658
rect 7593 69606 7605 69658
rect 7605 69606 7619 69658
rect 7643 69606 7657 69658
rect 7657 69606 7669 69658
rect 7669 69606 7699 69658
rect 7723 69606 7733 69658
rect 7733 69606 7779 69658
rect 7483 69604 7539 69606
rect 7563 69604 7619 69606
rect 7643 69604 7699 69606
rect 7723 69604 7779 69606
rect 5851 69114 5907 69116
rect 5931 69114 5987 69116
rect 6011 69114 6067 69116
rect 6091 69114 6147 69116
rect 5851 69062 5897 69114
rect 5897 69062 5907 69114
rect 5931 69062 5961 69114
rect 5961 69062 5973 69114
rect 5973 69062 5987 69114
rect 6011 69062 6025 69114
rect 6025 69062 6037 69114
rect 6037 69062 6067 69114
rect 6091 69062 6101 69114
rect 6101 69062 6147 69114
rect 5851 69060 5907 69062
rect 5931 69060 5987 69062
rect 6011 69060 6067 69062
rect 6091 69060 6147 69062
rect 5851 68026 5907 68028
rect 5931 68026 5987 68028
rect 6011 68026 6067 68028
rect 6091 68026 6147 68028
rect 5851 67974 5897 68026
rect 5897 67974 5907 68026
rect 5931 67974 5961 68026
rect 5961 67974 5973 68026
rect 5973 67974 5987 68026
rect 6011 67974 6025 68026
rect 6025 67974 6037 68026
rect 6037 67974 6067 68026
rect 6091 67974 6101 68026
rect 6101 67974 6147 68026
rect 5851 67972 5907 67974
rect 5931 67972 5987 67974
rect 6011 67972 6067 67974
rect 6091 67972 6147 67974
rect 5851 66938 5907 66940
rect 5931 66938 5987 66940
rect 6011 66938 6067 66940
rect 6091 66938 6147 66940
rect 5851 66886 5897 66938
rect 5897 66886 5907 66938
rect 5931 66886 5961 66938
rect 5961 66886 5973 66938
rect 5973 66886 5987 66938
rect 6011 66886 6025 66938
rect 6025 66886 6037 66938
rect 6037 66886 6067 66938
rect 6091 66886 6101 66938
rect 6101 66886 6147 66938
rect 5851 66884 5907 66886
rect 5931 66884 5987 66886
rect 6011 66884 6067 66886
rect 6091 66884 6147 66886
rect 5851 65850 5907 65852
rect 5931 65850 5987 65852
rect 6011 65850 6067 65852
rect 6091 65850 6147 65852
rect 5851 65798 5897 65850
rect 5897 65798 5907 65850
rect 5931 65798 5961 65850
rect 5961 65798 5973 65850
rect 5973 65798 5987 65850
rect 6011 65798 6025 65850
rect 6025 65798 6037 65850
rect 6037 65798 6067 65850
rect 6091 65798 6101 65850
rect 6101 65798 6147 65850
rect 5851 65796 5907 65798
rect 5931 65796 5987 65798
rect 6011 65796 6067 65798
rect 6091 65796 6147 65798
rect 5906 65628 5908 65648
rect 5908 65628 5960 65648
rect 5960 65628 5962 65648
rect 5906 65592 5962 65628
rect 5851 64762 5907 64764
rect 5931 64762 5987 64764
rect 6011 64762 6067 64764
rect 6091 64762 6147 64764
rect 5851 64710 5897 64762
rect 5897 64710 5907 64762
rect 5931 64710 5961 64762
rect 5961 64710 5973 64762
rect 5973 64710 5987 64762
rect 6011 64710 6025 64762
rect 6025 64710 6037 64762
rect 6037 64710 6067 64762
rect 6091 64710 6101 64762
rect 6101 64710 6147 64762
rect 5851 64708 5907 64710
rect 5931 64708 5987 64710
rect 6011 64708 6067 64710
rect 6091 64708 6147 64710
rect 5851 63674 5907 63676
rect 5931 63674 5987 63676
rect 6011 63674 6067 63676
rect 6091 63674 6147 63676
rect 5851 63622 5897 63674
rect 5897 63622 5907 63674
rect 5931 63622 5961 63674
rect 5961 63622 5973 63674
rect 5973 63622 5987 63674
rect 6011 63622 6025 63674
rect 6025 63622 6037 63674
rect 6037 63622 6067 63674
rect 6091 63622 6101 63674
rect 6101 63622 6147 63674
rect 5851 63620 5907 63622
rect 5931 63620 5987 63622
rect 6011 63620 6067 63622
rect 6091 63620 6147 63622
rect 5851 62586 5907 62588
rect 5931 62586 5987 62588
rect 6011 62586 6067 62588
rect 6091 62586 6147 62588
rect 5851 62534 5897 62586
rect 5897 62534 5907 62586
rect 5931 62534 5961 62586
rect 5961 62534 5973 62586
rect 5973 62534 5987 62586
rect 6011 62534 6025 62586
rect 6025 62534 6037 62586
rect 6037 62534 6067 62586
rect 6091 62534 6101 62586
rect 6101 62534 6147 62586
rect 5851 62532 5907 62534
rect 5931 62532 5987 62534
rect 6011 62532 6067 62534
rect 6091 62532 6147 62534
rect 5851 61498 5907 61500
rect 5931 61498 5987 61500
rect 6011 61498 6067 61500
rect 6091 61498 6147 61500
rect 5851 61446 5897 61498
rect 5897 61446 5907 61498
rect 5931 61446 5961 61498
rect 5961 61446 5973 61498
rect 5973 61446 5987 61498
rect 6011 61446 6025 61498
rect 6025 61446 6037 61498
rect 6037 61446 6067 61498
rect 6091 61446 6101 61498
rect 6101 61446 6147 61498
rect 5851 61444 5907 61446
rect 5931 61444 5987 61446
rect 6011 61444 6067 61446
rect 6091 61444 6147 61446
rect 5851 60410 5907 60412
rect 5931 60410 5987 60412
rect 6011 60410 6067 60412
rect 6091 60410 6147 60412
rect 5851 60358 5897 60410
rect 5897 60358 5907 60410
rect 5931 60358 5961 60410
rect 5961 60358 5973 60410
rect 5973 60358 5987 60410
rect 6011 60358 6025 60410
rect 6025 60358 6037 60410
rect 6037 60358 6067 60410
rect 6091 60358 6101 60410
rect 6101 60358 6147 60410
rect 5851 60356 5907 60358
rect 5931 60356 5987 60358
rect 6011 60356 6067 60358
rect 6091 60356 6147 60358
rect 5851 59322 5907 59324
rect 5931 59322 5987 59324
rect 6011 59322 6067 59324
rect 6091 59322 6147 59324
rect 5851 59270 5897 59322
rect 5897 59270 5907 59322
rect 5931 59270 5961 59322
rect 5961 59270 5973 59322
rect 5973 59270 5987 59322
rect 6011 59270 6025 59322
rect 6025 59270 6037 59322
rect 6037 59270 6067 59322
rect 6091 59270 6101 59322
rect 6101 59270 6147 59322
rect 5851 59268 5907 59270
rect 5931 59268 5987 59270
rect 6011 59268 6067 59270
rect 6091 59268 6147 59270
rect 5851 58234 5907 58236
rect 5931 58234 5987 58236
rect 6011 58234 6067 58236
rect 6091 58234 6147 58236
rect 5851 58182 5897 58234
rect 5897 58182 5907 58234
rect 5931 58182 5961 58234
rect 5961 58182 5973 58234
rect 5973 58182 5987 58234
rect 6011 58182 6025 58234
rect 6025 58182 6037 58234
rect 6037 58182 6067 58234
rect 6091 58182 6101 58234
rect 6101 58182 6147 58234
rect 5851 58180 5907 58182
rect 5931 58180 5987 58182
rect 6011 58180 6067 58182
rect 6091 58180 6147 58182
rect 5851 57146 5907 57148
rect 5931 57146 5987 57148
rect 6011 57146 6067 57148
rect 6091 57146 6147 57148
rect 5851 57094 5897 57146
rect 5897 57094 5907 57146
rect 5931 57094 5961 57146
rect 5961 57094 5973 57146
rect 5973 57094 5987 57146
rect 6011 57094 6025 57146
rect 6025 57094 6037 57146
rect 6037 57094 6067 57146
rect 6091 57094 6101 57146
rect 6101 57094 6147 57146
rect 5851 57092 5907 57094
rect 5931 57092 5987 57094
rect 6011 57092 6067 57094
rect 6091 57092 6147 57094
rect 5851 56058 5907 56060
rect 5931 56058 5987 56060
rect 6011 56058 6067 56060
rect 6091 56058 6147 56060
rect 5851 56006 5897 56058
rect 5897 56006 5907 56058
rect 5931 56006 5961 56058
rect 5961 56006 5973 56058
rect 5973 56006 5987 56058
rect 6011 56006 6025 56058
rect 6025 56006 6037 56058
rect 6037 56006 6067 56058
rect 6091 56006 6101 56058
rect 6101 56006 6147 56058
rect 5851 56004 5907 56006
rect 5931 56004 5987 56006
rect 6011 56004 6067 56006
rect 6091 56004 6147 56006
rect 5851 54970 5907 54972
rect 5931 54970 5987 54972
rect 6011 54970 6067 54972
rect 6091 54970 6147 54972
rect 5851 54918 5897 54970
rect 5897 54918 5907 54970
rect 5931 54918 5961 54970
rect 5961 54918 5973 54970
rect 5973 54918 5987 54970
rect 6011 54918 6025 54970
rect 6025 54918 6037 54970
rect 6037 54918 6067 54970
rect 6091 54918 6101 54970
rect 6101 54918 6147 54970
rect 5851 54916 5907 54918
rect 5931 54916 5987 54918
rect 6011 54916 6067 54918
rect 6091 54916 6147 54918
rect 5851 53882 5907 53884
rect 5931 53882 5987 53884
rect 6011 53882 6067 53884
rect 6091 53882 6147 53884
rect 5851 53830 5897 53882
rect 5897 53830 5907 53882
rect 5931 53830 5961 53882
rect 5961 53830 5973 53882
rect 5973 53830 5987 53882
rect 6011 53830 6025 53882
rect 6025 53830 6037 53882
rect 6037 53830 6067 53882
rect 6091 53830 6101 53882
rect 6101 53830 6147 53882
rect 5851 53828 5907 53830
rect 5931 53828 5987 53830
rect 6011 53828 6067 53830
rect 6091 53828 6147 53830
rect 5851 52794 5907 52796
rect 5931 52794 5987 52796
rect 6011 52794 6067 52796
rect 6091 52794 6147 52796
rect 5851 52742 5897 52794
rect 5897 52742 5907 52794
rect 5931 52742 5961 52794
rect 5961 52742 5973 52794
rect 5973 52742 5987 52794
rect 6011 52742 6025 52794
rect 6025 52742 6037 52794
rect 6037 52742 6067 52794
rect 6091 52742 6101 52794
rect 6101 52742 6147 52794
rect 5851 52740 5907 52742
rect 5931 52740 5987 52742
rect 6011 52740 6067 52742
rect 6091 52740 6147 52742
rect 5851 51706 5907 51708
rect 5931 51706 5987 51708
rect 6011 51706 6067 51708
rect 6091 51706 6147 51708
rect 5851 51654 5897 51706
rect 5897 51654 5907 51706
rect 5931 51654 5961 51706
rect 5961 51654 5973 51706
rect 5973 51654 5987 51706
rect 6011 51654 6025 51706
rect 6025 51654 6037 51706
rect 6037 51654 6067 51706
rect 6091 51654 6101 51706
rect 6101 51654 6147 51706
rect 5851 51652 5907 51654
rect 5931 51652 5987 51654
rect 6011 51652 6067 51654
rect 6091 51652 6147 51654
rect 5851 50618 5907 50620
rect 5931 50618 5987 50620
rect 6011 50618 6067 50620
rect 6091 50618 6147 50620
rect 5851 50566 5897 50618
rect 5897 50566 5907 50618
rect 5931 50566 5961 50618
rect 5961 50566 5973 50618
rect 5973 50566 5987 50618
rect 6011 50566 6025 50618
rect 6025 50566 6037 50618
rect 6037 50566 6067 50618
rect 6091 50566 6101 50618
rect 6101 50566 6147 50618
rect 5851 50564 5907 50566
rect 5931 50564 5987 50566
rect 6011 50564 6067 50566
rect 6091 50564 6147 50566
rect 5851 49530 5907 49532
rect 5931 49530 5987 49532
rect 6011 49530 6067 49532
rect 6091 49530 6147 49532
rect 5851 49478 5897 49530
rect 5897 49478 5907 49530
rect 5931 49478 5961 49530
rect 5961 49478 5973 49530
rect 5973 49478 5987 49530
rect 6011 49478 6025 49530
rect 6025 49478 6037 49530
rect 6037 49478 6067 49530
rect 6091 49478 6101 49530
rect 6101 49478 6147 49530
rect 5851 49476 5907 49478
rect 5931 49476 5987 49478
rect 6011 49476 6067 49478
rect 6091 49476 6147 49478
rect 5851 48442 5907 48444
rect 5931 48442 5987 48444
rect 6011 48442 6067 48444
rect 6091 48442 6147 48444
rect 5851 48390 5897 48442
rect 5897 48390 5907 48442
rect 5931 48390 5961 48442
rect 5961 48390 5973 48442
rect 5973 48390 5987 48442
rect 6011 48390 6025 48442
rect 6025 48390 6037 48442
rect 6037 48390 6067 48442
rect 6091 48390 6101 48442
rect 6101 48390 6147 48442
rect 5851 48388 5907 48390
rect 5931 48388 5987 48390
rect 6011 48388 6067 48390
rect 6091 48388 6147 48390
rect 5906 47504 5962 47560
rect 5851 47354 5907 47356
rect 5931 47354 5987 47356
rect 6011 47354 6067 47356
rect 6091 47354 6147 47356
rect 5851 47302 5897 47354
rect 5897 47302 5907 47354
rect 5931 47302 5961 47354
rect 5961 47302 5973 47354
rect 5973 47302 5987 47354
rect 6011 47302 6025 47354
rect 6025 47302 6037 47354
rect 6037 47302 6067 47354
rect 6091 47302 6101 47354
rect 6101 47302 6147 47354
rect 5851 47300 5907 47302
rect 5931 47300 5987 47302
rect 6011 47300 6067 47302
rect 6091 47300 6147 47302
rect 5851 46266 5907 46268
rect 5931 46266 5987 46268
rect 6011 46266 6067 46268
rect 6091 46266 6147 46268
rect 5851 46214 5897 46266
rect 5897 46214 5907 46266
rect 5931 46214 5961 46266
rect 5961 46214 5973 46266
rect 5973 46214 5987 46266
rect 6011 46214 6025 46266
rect 6025 46214 6037 46266
rect 6037 46214 6067 46266
rect 6091 46214 6101 46266
rect 6101 46214 6147 46266
rect 5851 46212 5907 46214
rect 5931 46212 5987 46214
rect 6011 46212 6067 46214
rect 6091 46212 6147 46214
rect 5851 45178 5907 45180
rect 5931 45178 5987 45180
rect 6011 45178 6067 45180
rect 6091 45178 6147 45180
rect 5851 45126 5897 45178
rect 5897 45126 5907 45178
rect 5931 45126 5961 45178
rect 5961 45126 5973 45178
rect 5973 45126 5987 45178
rect 6011 45126 6025 45178
rect 6025 45126 6037 45178
rect 6037 45126 6067 45178
rect 6091 45126 6101 45178
rect 6101 45126 6147 45178
rect 5851 45124 5907 45126
rect 5931 45124 5987 45126
rect 6011 45124 6067 45126
rect 6091 45124 6147 45126
rect 5851 44090 5907 44092
rect 5931 44090 5987 44092
rect 6011 44090 6067 44092
rect 6091 44090 6147 44092
rect 5851 44038 5897 44090
rect 5897 44038 5907 44090
rect 5931 44038 5961 44090
rect 5961 44038 5973 44090
rect 5973 44038 5987 44090
rect 6011 44038 6025 44090
rect 6025 44038 6037 44090
rect 6037 44038 6067 44090
rect 6091 44038 6101 44090
rect 6101 44038 6147 44090
rect 5851 44036 5907 44038
rect 5931 44036 5987 44038
rect 6011 44036 6067 44038
rect 6091 44036 6147 44038
rect 5851 43002 5907 43004
rect 5931 43002 5987 43004
rect 6011 43002 6067 43004
rect 6091 43002 6147 43004
rect 5851 42950 5897 43002
rect 5897 42950 5907 43002
rect 5931 42950 5961 43002
rect 5961 42950 5973 43002
rect 5973 42950 5987 43002
rect 6011 42950 6025 43002
rect 6025 42950 6037 43002
rect 6037 42950 6067 43002
rect 6091 42950 6101 43002
rect 6101 42950 6147 43002
rect 5851 42948 5907 42950
rect 5931 42948 5987 42950
rect 6011 42948 6067 42950
rect 6091 42948 6147 42950
rect 5851 41914 5907 41916
rect 5931 41914 5987 41916
rect 6011 41914 6067 41916
rect 6091 41914 6147 41916
rect 5851 41862 5897 41914
rect 5897 41862 5907 41914
rect 5931 41862 5961 41914
rect 5961 41862 5973 41914
rect 5973 41862 5987 41914
rect 6011 41862 6025 41914
rect 6025 41862 6037 41914
rect 6037 41862 6067 41914
rect 6091 41862 6101 41914
rect 6101 41862 6147 41914
rect 5851 41860 5907 41862
rect 5931 41860 5987 41862
rect 6011 41860 6067 41862
rect 6091 41860 6147 41862
rect 5851 40826 5907 40828
rect 5931 40826 5987 40828
rect 6011 40826 6067 40828
rect 6091 40826 6147 40828
rect 5851 40774 5897 40826
rect 5897 40774 5907 40826
rect 5931 40774 5961 40826
rect 5961 40774 5973 40826
rect 5973 40774 5987 40826
rect 6011 40774 6025 40826
rect 6025 40774 6037 40826
rect 6037 40774 6067 40826
rect 6091 40774 6101 40826
rect 6101 40774 6147 40826
rect 5851 40772 5907 40774
rect 5931 40772 5987 40774
rect 6011 40772 6067 40774
rect 6091 40772 6147 40774
rect 5851 39738 5907 39740
rect 5931 39738 5987 39740
rect 6011 39738 6067 39740
rect 6091 39738 6147 39740
rect 5851 39686 5897 39738
rect 5897 39686 5907 39738
rect 5931 39686 5961 39738
rect 5961 39686 5973 39738
rect 5973 39686 5987 39738
rect 6011 39686 6025 39738
rect 6025 39686 6037 39738
rect 6037 39686 6067 39738
rect 6091 39686 6101 39738
rect 6101 39686 6147 39738
rect 5851 39684 5907 39686
rect 5931 39684 5987 39686
rect 6011 39684 6067 39686
rect 6091 39684 6147 39686
rect 5851 38650 5907 38652
rect 5931 38650 5987 38652
rect 6011 38650 6067 38652
rect 6091 38650 6147 38652
rect 5851 38598 5897 38650
rect 5897 38598 5907 38650
rect 5931 38598 5961 38650
rect 5961 38598 5973 38650
rect 5973 38598 5987 38650
rect 6011 38598 6025 38650
rect 6025 38598 6037 38650
rect 6037 38598 6067 38650
rect 6091 38598 6101 38650
rect 6101 38598 6147 38650
rect 5851 38596 5907 38598
rect 5931 38596 5987 38598
rect 6011 38596 6067 38598
rect 6091 38596 6147 38598
rect 5851 37562 5907 37564
rect 5931 37562 5987 37564
rect 6011 37562 6067 37564
rect 6091 37562 6147 37564
rect 5851 37510 5897 37562
rect 5897 37510 5907 37562
rect 5931 37510 5961 37562
rect 5961 37510 5973 37562
rect 5973 37510 5987 37562
rect 6011 37510 6025 37562
rect 6025 37510 6037 37562
rect 6037 37510 6067 37562
rect 6091 37510 6101 37562
rect 6101 37510 6147 37562
rect 5851 37508 5907 37510
rect 5931 37508 5987 37510
rect 6011 37508 6067 37510
rect 6091 37508 6147 37510
rect 5851 36474 5907 36476
rect 5931 36474 5987 36476
rect 6011 36474 6067 36476
rect 6091 36474 6147 36476
rect 5851 36422 5897 36474
rect 5897 36422 5907 36474
rect 5931 36422 5961 36474
rect 5961 36422 5973 36474
rect 5973 36422 5987 36474
rect 6011 36422 6025 36474
rect 6025 36422 6037 36474
rect 6037 36422 6067 36474
rect 6091 36422 6101 36474
rect 6101 36422 6147 36474
rect 5851 36420 5907 36422
rect 5931 36420 5987 36422
rect 6011 36420 6067 36422
rect 6091 36420 6147 36422
rect 5851 35386 5907 35388
rect 5931 35386 5987 35388
rect 6011 35386 6067 35388
rect 6091 35386 6147 35388
rect 5851 35334 5897 35386
rect 5897 35334 5907 35386
rect 5931 35334 5961 35386
rect 5961 35334 5973 35386
rect 5973 35334 5987 35386
rect 6011 35334 6025 35386
rect 6025 35334 6037 35386
rect 6037 35334 6067 35386
rect 6091 35334 6101 35386
rect 6101 35334 6147 35386
rect 5851 35332 5907 35334
rect 5931 35332 5987 35334
rect 6011 35332 6067 35334
rect 6091 35332 6147 35334
rect 5851 34298 5907 34300
rect 5931 34298 5987 34300
rect 6011 34298 6067 34300
rect 6091 34298 6147 34300
rect 5851 34246 5897 34298
rect 5897 34246 5907 34298
rect 5931 34246 5961 34298
rect 5961 34246 5973 34298
rect 5973 34246 5987 34298
rect 6011 34246 6025 34298
rect 6025 34246 6037 34298
rect 6037 34246 6067 34298
rect 6091 34246 6101 34298
rect 6101 34246 6147 34298
rect 5851 34244 5907 34246
rect 5931 34244 5987 34246
rect 6011 34244 6067 34246
rect 6091 34244 6147 34246
rect 5851 33210 5907 33212
rect 5931 33210 5987 33212
rect 6011 33210 6067 33212
rect 6091 33210 6147 33212
rect 5851 33158 5897 33210
rect 5897 33158 5907 33210
rect 5931 33158 5961 33210
rect 5961 33158 5973 33210
rect 5973 33158 5987 33210
rect 6011 33158 6025 33210
rect 6025 33158 6037 33210
rect 6037 33158 6067 33210
rect 6091 33158 6101 33210
rect 6101 33158 6147 33210
rect 5851 33156 5907 33158
rect 5931 33156 5987 33158
rect 6011 33156 6067 33158
rect 6091 33156 6147 33158
rect 5851 32122 5907 32124
rect 5931 32122 5987 32124
rect 6011 32122 6067 32124
rect 6091 32122 6147 32124
rect 5851 32070 5897 32122
rect 5897 32070 5907 32122
rect 5931 32070 5961 32122
rect 5961 32070 5973 32122
rect 5973 32070 5987 32122
rect 6011 32070 6025 32122
rect 6025 32070 6037 32122
rect 6037 32070 6067 32122
rect 6091 32070 6101 32122
rect 6101 32070 6147 32122
rect 5851 32068 5907 32070
rect 5931 32068 5987 32070
rect 6011 32068 6067 32070
rect 6091 32068 6147 32070
rect 5851 31034 5907 31036
rect 5931 31034 5987 31036
rect 6011 31034 6067 31036
rect 6091 31034 6147 31036
rect 5851 30982 5897 31034
rect 5897 30982 5907 31034
rect 5931 30982 5961 31034
rect 5961 30982 5973 31034
rect 5973 30982 5987 31034
rect 6011 30982 6025 31034
rect 6025 30982 6037 31034
rect 6037 30982 6067 31034
rect 6091 30982 6101 31034
rect 6101 30982 6147 31034
rect 5851 30980 5907 30982
rect 5931 30980 5987 30982
rect 6011 30980 6067 30982
rect 6091 30980 6147 30982
rect 5851 29946 5907 29948
rect 5931 29946 5987 29948
rect 6011 29946 6067 29948
rect 6091 29946 6147 29948
rect 5851 29894 5897 29946
rect 5897 29894 5907 29946
rect 5931 29894 5961 29946
rect 5961 29894 5973 29946
rect 5973 29894 5987 29946
rect 6011 29894 6025 29946
rect 6025 29894 6037 29946
rect 6037 29894 6067 29946
rect 6091 29894 6101 29946
rect 6101 29894 6147 29946
rect 5851 29892 5907 29894
rect 5931 29892 5987 29894
rect 6011 29892 6067 29894
rect 6091 29892 6147 29894
rect 5851 28858 5907 28860
rect 5931 28858 5987 28860
rect 6011 28858 6067 28860
rect 6091 28858 6147 28860
rect 5851 28806 5897 28858
rect 5897 28806 5907 28858
rect 5931 28806 5961 28858
rect 5961 28806 5973 28858
rect 5973 28806 5987 28858
rect 6011 28806 6025 28858
rect 6025 28806 6037 28858
rect 6037 28806 6067 28858
rect 6091 28806 6101 28858
rect 6101 28806 6147 28858
rect 5851 28804 5907 28806
rect 5931 28804 5987 28806
rect 6011 28804 6067 28806
rect 6091 28804 6147 28806
rect 5851 27770 5907 27772
rect 5931 27770 5987 27772
rect 6011 27770 6067 27772
rect 6091 27770 6147 27772
rect 5851 27718 5897 27770
rect 5897 27718 5907 27770
rect 5931 27718 5961 27770
rect 5961 27718 5973 27770
rect 5973 27718 5987 27770
rect 6011 27718 6025 27770
rect 6025 27718 6037 27770
rect 6037 27718 6067 27770
rect 6091 27718 6101 27770
rect 6101 27718 6147 27770
rect 5851 27716 5907 27718
rect 5931 27716 5987 27718
rect 6011 27716 6067 27718
rect 6091 27716 6147 27718
rect 5851 26682 5907 26684
rect 5931 26682 5987 26684
rect 6011 26682 6067 26684
rect 6091 26682 6147 26684
rect 5851 26630 5897 26682
rect 5897 26630 5907 26682
rect 5931 26630 5961 26682
rect 5961 26630 5973 26682
rect 5973 26630 5987 26682
rect 6011 26630 6025 26682
rect 6025 26630 6037 26682
rect 6037 26630 6067 26682
rect 6091 26630 6101 26682
rect 6101 26630 6147 26682
rect 5851 26628 5907 26630
rect 5931 26628 5987 26630
rect 6011 26628 6067 26630
rect 6091 26628 6147 26630
rect 5851 25594 5907 25596
rect 5931 25594 5987 25596
rect 6011 25594 6067 25596
rect 6091 25594 6147 25596
rect 5851 25542 5897 25594
rect 5897 25542 5907 25594
rect 5931 25542 5961 25594
rect 5961 25542 5973 25594
rect 5973 25542 5987 25594
rect 6011 25542 6025 25594
rect 6025 25542 6037 25594
rect 6037 25542 6067 25594
rect 6091 25542 6101 25594
rect 6101 25542 6147 25594
rect 5851 25540 5907 25542
rect 5931 25540 5987 25542
rect 6011 25540 6067 25542
rect 6091 25540 6147 25542
rect 5851 24506 5907 24508
rect 5931 24506 5987 24508
rect 6011 24506 6067 24508
rect 6091 24506 6147 24508
rect 5851 24454 5897 24506
rect 5897 24454 5907 24506
rect 5931 24454 5961 24506
rect 5961 24454 5973 24506
rect 5973 24454 5987 24506
rect 6011 24454 6025 24506
rect 6025 24454 6037 24506
rect 6037 24454 6067 24506
rect 6091 24454 6101 24506
rect 6101 24454 6147 24506
rect 5851 24452 5907 24454
rect 5931 24452 5987 24454
rect 6011 24452 6067 24454
rect 6091 24452 6147 24454
rect 5851 23418 5907 23420
rect 5931 23418 5987 23420
rect 6011 23418 6067 23420
rect 6091 23418 6147 23420
rect 5851 23366 5897 23418
rect 5897 23366 5907 23418
rect 5931 23366 5961 23418
rect 5961 23366 5973 23418
rect 5973 23366 5987 23418
rect 6011 23366 6025 23418
rect 6025 23366 6037 23418
rect 6037 23366 6067 23418
rect 6091 23366 6101 23418
rect 6101 23366 6147 23418
rect 5851 23364 5907 23366
rect 5931 23364 5987 23366
rect 6011 23364 6067 23366
rect 6091 23364 6147 23366
rect 5851 22330 5907 22332
rect 5931 22330 5987 22332
rect 6011 22330 6067 22332
rect 6091 22330 6147 22332
rect 5851 22278 5897 22330
rect 5897 22278 5907 22330
rect 5931 22278 5961 22330
rect 5961 22278 5973 22330
rect 5973 22278 5987 22330
rect 6011 22278 6025 22330
rect 6025 22278 6037 22330
rect 6037 22278 6067 22330
rect 6091 22278 6101 22330
rect 6101 22278 6147 22330
rect 5851 22276 5907 22278
rect 5931 22276 5987 22278
rect 6011 22276 6067 22278
rect 6091 22276 6147 22278
rect 5851 21242 5907 21244
rect 5931 21242 5987 21244
rect 6011 21242 6067 21244
rect 6091 21242 6147 21244
rect 5851 21190 5897 21242
rect 5897 21190 5907 21242
rect 5931 21190 5961 21242
rect 5961 21190 5973 21242
rect 5973 21190 5987 21242
rect 6011 21190 6025 21242
rect 6025 21190 6037 21242
rect 6037 21190 6067 21242
rect 6091 21190 6101 21242
rect 6101 21190 6147 21242
rect 5851 21188 5907 21190
rect 5931 21188 5987 21190
rect 6011 21188 6067 21190
rect 6091 21188 6147 21190
rect 5851 20154 5907 20156
rect 5931 20154 5987 20156
rect 6011 20154 6067 20156
rect 6091 20154 6147 20156
rect 5851 20102 5897 20154
rect 5897 20102 5907 20154
rect 5931 20102 5961 20154
rect 5961 20102 5973 20154
rect 5973 20102 5987 20154
rect 6011 20102 6025 20154
rect 6025 20102 6037 20154
rect 6037 20102 6067 20154
rect 6091 20102 6101 20154
rect 6101 20102 6147 20154
rect 5851 20100 5907 20102
rect 5931 20100 5987 20102
rect 6011 20100 6067 20102
rect 6091 20100 6147 20102
rect 5851 19066 5907 19068
rect 5931 19066 5987 19068
rect 6011 19066 6067 19068
rect 6091 19066 6147 19068
rect 5851 19014 5897 19066
rect 5897 19014 5907 19066
rect 5931 19014 5961 19066
rect 5961 19014 5973 19066
rect 5973 19014 5987 19066
rect 6011 19014 6025 19066
rect 6025 19014 6037 19066
rect 6037 19014 6067 19066
rect 6091 19014 6101 19066
rect 6101 19014 6147 19066
rect 5851 19012 5907 19014
rect 5931 19012 5987 19014
rect 6011 19012 6067 19014
rect 6091 19012 6147 19014
rect 5851 17978 5907 17980
rect 5931 17978 5987 17980
rect 6011 17978 6067 17980
rect 6091 17978 6147 17980
rect 5851 17926 5897 17978
rect 5897 17926 5907 17978
rect 5931 17926 5961 17978
rect 5961 17926 5973 17978
rect 5973 17926 5987 17978
rect 6011 17926 6025 17978
rect 6025 17926 6037 17978
rect 6037 17926 6067 17978
rect 6091 17926 6101 17978
rect 6101 17926 6147 17978
rect 5851 17924 5907 17926
rect 5931 17924 5987 17926
rect 6011 17924 6067 17926
rect 6091 17924 6147 17926
rect 5851 16890 5907 16892
rect 5931 16890 5987 16892
rect 6011 16890 6067 16892
rect 6091 16890 6147 16892
rect 5851 16838 5897 16890
rect 5897 16838 5907 16890
rect 5931 16838 5961 16890
rect 5961 16838 5973 16890
rect 5973 16838 5987 16890
rect 6011 16838 6025 16890
rect 6025 16838 6037 16890
rect 6037 16838 6067 16890
rect 6091 16838 6101 16890
rect 6101 16838 6147 16890
rect 5851 16836 5907 16838
rect 5931 16836 5987 16838
rect 6011 16836 6067 16838
rect 6091 16836 6147 16838
rect 5851 15802 5907 15804
rect 5931 15802 5987 15804
rect 6011 15802 6067 15804
rect 6091 15802 6147 15804
rect 5851 15750 5897 15802
rect 5897 15750 5907 15802
rect 5931 15750 5961 15802
rect 5961 15750 5973 15802
rect 5973 15750 5987 15802
rect 6011 15750 6025 15802
rect 6025 15750 6037 15802
rect 6037 15750 6067 15802
rect 6091 15750 6101 15802
rect 6101 15750 6147 15802
rect 5851 15748 5907 15750
rect 5931 15748 5987 15750
rect 6011 15748 6067 15750
rect 6091 15748 6147 15750
rect 5851 14714 5907 14716
rect 5931 14714 5987 14716
rect 6011 14714 6067 14716
rect 6091 14714 6147 14716
rect 5851 14662 5897 14714
rect 5897 14662 5907 14714
rect 5931 14662 5961 14714
rect 5961 14662 5973 14714
rect 5973 14662 5987 14714
rect 6011 14662 6025 14714
rect 6025 14662 6037 14714
rect 6037 14662 6067 14714
rect 6091 14662 6101 14714
rect 6101 14662 6147 14714
rect 5851 14660 5907 14662
rect 5931 14660 5987 14662
rect 6011 14660 6067 14662
rect 6091 14660 6147 14662
rect 5851 13626 5907 13628
rect 5931 13626 5987 13628
rect 6011 13626 6067 13628
rect 6091 13626 6147 13628
rect 5851 13574 5897 13626
rect 5897 13574 5907 13626
rect 5931 13574 5961 13626
rect 5961 13574 5973 13626
rect 5973 13574 5987 13626
rect 6011 13574 6025 13626
rect 6025 13574 6037 13626
rect 6037 13574 6067 13626
rect 6091 13574 6101 13626
rect 6101 13574 6147 13626
rect 5851 13572 5907 13574
rect 5931 13572 5987 13574
rect 6011 13572 6067 13574
rect 6091 13572 6147 13574
rect 5851 12538 5907 12540
rect 5931 12538 5987 12540
rect 6011 12538 6067 12540
rect 6091 12538 6147 12540
rect 5851 12486 5897 12538
rect 5897 12486 5907 12538
rect 5931 12486 5961 12538
rect 5961 12486 5973 12538
rect 5973 12486 5987 12538
rect 6011 12486 6025 12538
rect 6025 12486 6037 12538
rect 6037 12486 6067 12538
rect 6091 12486 6101 12538
rect 6101 12486 6147 12538
rect 5851 12484 5907 12486
rect 5931 12484 5987 12486
rect 6011 12484 6067 12486
rect 6091 12484 6147 12486
rect 5851 11450 5907 11452
rect 5931 11450 5987 11452
rect 6011 11450 6067 11452
rect 6091 11450 6147 11452
rect 5851 11398 5897 11450
rect 5897 11398 5907 11450
rect 5931 11398 5961 11450
rect 5961 11398 5973 11450
rect 5973 11398 5987 11450
rect 6011 11398 6025 11450
rect 6025 11398 6037 11450
rect 6037 11398 6067 11450
rect 6091 11398 6101 11450
rect 6101 11398 6147 11450
rect 5851 11396 5907 11398
rect 5931 11396 5987 11398
rect 6011 11396 6067 11398
rect 6091 11396 6147 11398
rect 5851 10362 5907 10364
rect 5931 10362 5987 10364
rect 6011 10362 6067 10364
rect 6091 10362 6147 10364
rect 5851 10310 5897 10362
rect 5897 10310 5907 10362
rect 5931 10310 5961 10362
rect 5961 10310 5973 10362
rect 5973 10310 5987 10362
rect 6011 10310 6025 10362
rect 6025 10310 6037 10362
rect 6037 10310 6067 10362
rect 6091 10310 6101 10362
rect 6101 10310 6147 10362
rect 5851 10308 5907 10310
rect 5931 10308 5987 10310
rect 6011 10308 6067 10310
rect 6091 10308 6147 10310
rect 5851 9274 5907 9276
rect 5931 9274 5987 9276
rect 6011 9274 6067 9276
rect 6091 9274 6147 9276
rect 5851 9222 5897 9274
rect 5897 9222 5907 9274
rect 5931 9222 5961 9274
rect 5961 9222 5973 9274
rect 5973 9222 5987 9274
rect 6011 9222 6025 9274
rect 6025 9222 6037 9274
rect 6037 9222 6067 9274
rect 6091 9222 6101 9274
rect 6101 9222 6147 9274
rect 5851 9220 5907 9222
rect 5931 9220 5987 9222
rect 6011 9220 6067 9222
rect 6091 9220 6147 9222
rect 6734 43696 6790 43752
rect 7483 68570 7539 68572
rect 7563 68570 7619 68572
rect 7643 68570 7699 68572
rect 7723 68570 7779 68572
rect 7483 68518 7529 68570
rect 7529 68518 7539 68570
rect 7563 68518 7593 68570
rect 7593 68518 7605 68570
rect 7605 68518 7619 68570
rect 7643 68518 7657 68570
rect 7657 68518 7669 68570
rect 7669 68518 7699 68570
rect 7723 68518 7733 68570
rect 7733 68518 7779 68570
rect 7483 68516 7539 68518
rect 7563 68516 7619 68518
rect 7643 68516 7699 68518
rect 7723 68516 7779 68518
rect 7483 67482 7539 67484
rect 7563 67482 7619 67484
rect 7643 67482 7699 67484
rect 7723 67482 7779 67484
rect 7483 67430 7529 67482
rect 7529 67430 7539 67482
rect 7563 67430 7593 67482
rect 7593 67430 7605 67482
rect 7605 67430 7619 67482
rect 7643 67430 7657 67482
rect 7657 67430 7669 67482
rect 7669 67430 7699 67482
rect 7723 67430 7733 67482
rect 7733 67430 7779 67482
rect 7483 67428 7539 67430
rect 7563 67428 7619 67430
rect 7643 67428 7699 67430
rect 7723 67428 7779 67430
rect 7483 66394 7539 66396
rect 7563 66394 7619 66396
rect 7643 66394 7699 66396
rect 7723 66394 7779 66396
rect 7483 66342 7529 66394
rect 7529 66342 7539 66394
rect 7563 66342 7593 66394
rect 7593 66342 7605 66394
rect 7605 66342 7619 66394
rect 7643 66342 7657 66394
rect 7657 66342 7669 66394
rect 7669 66342 7699 66394
rect 7723 66342 7733 66394
rect 7733 66342 7779 66394
rect 7483 66340 7539 66342
rect 7563 66340 7619 66342
rect 7643 66340 7699 66342
rect 7723 66340 7779 66342
rect 7194 66136 7250 66192
rect 7483 65306 7539 65308
rect 7563 65306 7619 65308
rect 7643 65306 7699 65308
rect 7723 65306 7779 65308
rect 7483 65254 7529 65306
rect 7529 65254 7539 65306
rect 7563 65254 7593 65306
rect 7593 65254 7605 65306
rect 7605 65254 7619 65306
rect 7643 65254 7657 65306
rect 7657 65254 7669 65306
rect 7669 65254 7699 65306
rect 7723 65254 7733 65306
rect 7733 65254 7779 65306
rect 7483 65252 7539 65254
rect 7563 65252 7619 65254
rect 7643 65252 7699 65254
rect 7723 65252 7779 65254
rect 7483 64218 7539 64220
rect 7563 64218 7619 64220
rect 7643 64218 7699 64220
rect 7723 64218 7779 64220
rect 7483 64166 7529 64218
rect 7529 64166 7539 64218
rect 7563 64166 7593 64218
rect 7593 64166 7605 64218
rect 7605 64166 7619 64218
rect 7643 64166 7657 64218
rect 7657 64166 7669 64218
rect 7669 64166 7699 64218
rect 7723 64166 7733 64218
rect 7733 64166 7779 64218
rect 7483 64164 7539 64166
rect 7563 64164 7619 64166
rect 7643 64164 7699 64166
rect 7723 64164 7779 64166
rect 7483 63130 7539 63132
rect 7563 63130 7619 63132
rect 7643 63130 7699 63132
rect 7723 63130 7779 63132
rect 7483 63078 7529 63130
rect 7529 63078 7539 63130
rect 7563 63078 7593 63130
rect 7593 63078 7605 63130
rect 7605 63078 7619 63130
rect 7643 63078 7657 63130
rect 7657 63078 7669 63130
rect 7669 63078 7699 63130
rect 7723 63078 7733 63130
rect 7733 63078 7779 63130
rect 7483 63076 7539 63078
rect 7563 63076 7619 63078
rect 7643 63076 7699 63078
rect 7723 63076 7779 63078
rect 7483 62042 7539 62044
rect 7563 62042 7619 62044
rect 7643 62042 7699 62044
rect 7723 62042 7779 62044
rect 7483 61990 7529 62042
rect 7529 61990 7539 62042
rect 7563 61990 7593 62042
rect 7593 61990 7605 62042
rect 7605 61990 7619 62042
rect 7643 61990 7657 62042
rect 7657 61990 7669 62042
rect 7669 61990 7699 62042
rect 7723 61990 7733 62042
rect 7733 61990 7779 62042
rect 7483 61988 7539 61990
rect 7563 61988 7619 61990
rect 7643 61988 7699 61990
rect 7723 61988 7779 61990
rect 7483 60954 7539 60956
rect 7563 60954 7619 60956
rect 7643 60954 7699 60956
rect 7723 60954 7779 60956
rect 7483 60902 7529 60954
rect 7529 60902 7539 60954
rect 7563 60902 7593 60954
rect 7593 60902 7605 60954
rect 7605 60902 7619 60954
rect 7643 60902 7657 60954
rect 7657 60902 7669 60954
rect 7669 60902 7699 60954
rect 7723 60902 7733 60954
rect 7733 60902 7779 60954
rect 7483 60900 7539 60902
rect 7563 60900 7619 60902
rect 7643 60900 7699 60902
rect 7723 60900 7779 60902
rect 7483 59866 7539 59868
rect 7563 59866 7619 59868
rect 7643 59866 7699 59868
rect 7723 59866 7779 59868
rect 7483 59814 7529 59866
rect 7529 59814 7539 59866
rect 7563 59814 7593 59866
rect 7593 59814 7605 59866
rect 7605 59814 7619 59866
rect 7643 59814 7657 59866
rect 7657 59814 7669 59866
rect 7669 59814 7699 59866
rect 7723 59814 7733 59866
rect 7733 59814 7779 59866
rect 7483 59812 7539 59814
rect 7563 59812 7619 59814
rect 7643 59812 7699 59814
rect 7723 59812 7779 59814
rect 7483 58778 7539 58780
rect 7563 58778 7619 58780
rect 7643 58778 7699 58780
rect 7723 58778 7779 58780
rect 7483 58726 7529 58778
rect 7529 58726 7539 58778
rect 7563 58726 7593 58778
rect 7593 58726 7605 58778
rect 7605 58726 7619 58778
rect 7643 58726 7657 58778
rect 7657 58726 7669 58778
rect 7669 58726 7699 58778
rect 7723 58726 7733 58778
rect 7733 58726 7779 58778
rect 7483 58724 7539 58726
rect 7563 58724 7619 58726
rect 7643 58724 7699 58726
rect 7723 58724 7779 58726
rect 7483 57690 7539 57692
rect 7563 57690 7619 57692
rect 7643 57690 7699 57692
rect 7723 57690 7779 57692
rect 7483 57638 7529 57690
rect 7529 57638 7539 57690
rect 7563 57638 7593 57690
rect 7593 57638 7605 57690
rect 7605 57638 7619 57690
rect 7643 57638 7657 57690
rect 7657 57638 7669 57690
rect 7669 57638 7699 57690
rect 7723 57638 7733 57690
rect 7733 57638 7779 57690
rect 7483 57636 7539 57638
rect 7563 57636 7619 57638
rect 7643 57636 7699 57638
rect 7723 57636 7779 57638
rect 7483 56602 7539 56604
rect 7563 56602 7619 56604
rect 7643 56602 7699 56604
rect 7723 56602 7779 56604
rect 7483 56550 7529 56602
rect 7529 56550 7539 56602
rect 7563 56550 7593 56602
rect 7593 56550 7605 56602
rect 7605 56550 7619 56602
rect 7643 56550 7657 56602
rect 7657 56550 7669 56602
rect 7669 56550 7699 56602
rect 7723 56550 7733 56602
rect 7733 56550 7779 56602
rect 7483 56548 7539 56550
rect 7563 56548 7619 56550
rect 7643 56548 7699 56550
rect 7723 56548 7779 56550
rect 7483 55514 7539 55516
rect 7563 55514 7619 55516
rect 7643 55514 7699 55516
rect 7723 55514 7779 55516
rect 7483 55462 7529 55514
rect 7529 55462 7539 55514
rect 7563 55462 7593 55514
rect 7593 55462 7605 55514
rect 7605 55462 7619 55514
rect 7643 55462 7657 55514
rect 7657 55462 7669 55514
rect 7669 55462 7699 55514
rect 7723 55462 7733 55514
rect 7733 55462 7779 55514
rect 7483 55460 7539 55462
rect 7563 55460 7619 55462
rect 7643 55460 7699 55462
rect 7723 55460 7779 55462
rect 7483 54426 7539 54428
rect 7563 54426 7619 54428
rect 7643 54426 7699 54428
rect 7723 54426 7779 54428
rect 7483 54374 7529 54426
rect 7529 54374 7539 54426
rect 7563 54374 7593 54426
rect 7593 54374 7605 54426
rect 7605 54374 7619 54426
rect 7643 54374 7657 54426
rect 7657 54374 7669 54426
rect 7669 54374 7699 54426
rect 7723 54374 7733 54426
rect 7733 54374 7779 54426
rect 7483 54372 7539 54374
rect 7563 54372 7619 54374
rect 7643 54372 7699 54374
rect 7723 54372 7779 54374
rect 7483 53338 7539 53340
rect 7563 53338 7619 53340
rect 7643 53338 7699 53340
rect 7723 53338 7779 53340
rect 7483 53286 7529 53338
rect 7529 53286 7539 53338
rect 7563 53286 7593 53338
rect 7593 53286 7605 53338
rect 7605 53286 7619 53338
rect 7643 53286 7657 53338
rect 7657 53286 7669 53338
rect 7669 53286 7699 53338
rect 7723 53286 7733 53338
rect 7733 53286 7779 53338
rect 7483 53284 7539 53286
rect 7563 53284 7619 53286
rect 7643 53284 7699 53286
rect 7723 53284 7779 53286
rect 7483 52250 7539 52252
rect 7563 52250 7619 52252
rect 7643 52250 7699 52252
rect 7723 52250 7779 52252
rect 7483 52198 7529 52250
rect 7529 52198 7539 52250
rect 7563 52198 7593 52250
rect 7593 52198 7605 52250
rect 7605 52198 7619 52250
rect 7643 52198 7657 52250
rect 7657 52198 7669 52250
rect 7669 52198 7699 52250
rect 7723 52198 7733 52250
rect 7733 52198 7779 52250
rect 7483 52196 7539 52198
rect 7563 52196 7619 52198
rect 7643 52196 7699 52198
rect 7723 52196 7779 52198
rect 7483 51162 7539 51164
rect 7563 51162 7619 51164
rect 7643 51162 7699 51164
rect 7723 51162 7779 51164
rect 7483 51110 7529 51162
rect 7529 51110 7539 51162
rect 7563 51110 7593 51162
rect 7593 51110 7605 51162
rect 7605 51110 7619 51162
rect 7643 51110 7657 51162
rect 7657 51110 7669 51162
rect 7669 51110 7699 51162
rect 7723 51110 7733 51162
rect 7733 51110 7779 51162
rect 7483 51108 7539 51110
rect 7563 51108 7619 51110
rect 7643 51108 7699 51110
rect 7723 51108 7779 51110
rect 7483 50074 7539 50076
rect 7563 50074 7619 50076
rect 7643 50074 7699 50076
rect 7723 50074 7779 50076
rect 7483 50022 7529 50074
rect 7529 50022 7539 50074
rect 7563 50022 7593 50074
rect 7593 50022 7605 50074
rect 7605 50022 7619 50074
rect 7643 50022 7657 50074
rect 7657 50022 7669 50074
rect 7669 50022 7699 50074
rect 7723 50022 7733 50074
rect 7733 50022 7779 50074
rect 7483 50020 7539 50022
rect 7563 50020 7619 50022
rect 7643 50020 7699 50022
rect 7723 50020 7779 50022
rect 7483 48986 7539 48988
rect 7563 48986 7619 48988
rect 7643 48986 7699 48988
rect 7723 48986 7779 48988
rect 7483 48934 7529 48986
rect 7529 48934 7539 48986
rect 7563 48934 7593 48986
rect 7593 48934 7605 48986
rect 7605 48934 7619 48986
rect 7643 48934 7657 48986
rect 7657 48934 7669 48986
rect 7669 48934 7699 48986
rect 7723 48934 7733 48986
rect 7733 48934 7779 48986
rect 7483 48932 7539 48934
rect 7563 48932 7619 48934
rect 7643 48932 7699 48934
rect 7723 48932 7779 48934
rect 7483 47898 7539 47900
rect 7563 47898 7619 47900
rect 7643 47898 7699 47900
rect 7723 47898 7779 47900
rect 7483 47846 7529 47898
rect 7529 47846 7539 47898
rect 7563 47846 7593 47898
rect 7593 47846 7605 47898
rect 7605 47846 7619 47898
rect 7643 47846 7657 47898
rect 7657 47846 7669 47898
rect 7669 47846 7699 47898
rect 7723 47846 7733 47898
rect 7733 47846 7779 47898
rect 7483 47844 7539 47846
rect 7563 47844 7619 47846
rect 7643 47844 7699 47846
rect 7723 47844 7779 47846
rect 7483 46810 7539 46812
rect 7563 46810 7619 46812
rect 7643 46810 7699 46812
rect 7723 46810 7779 46812
rect 7483 46758 7529 46810
rect 7529 46758 7539 46810
rect 7563 46758 7593 46810
rect 7593 46758 7605 46810
rect 7605 46758 7619 46810
rect 7643 46758 7657 46810
rect 7657 46758 7669 46810
rect 7669 46758 7699 46810
rect 7723 46758 7733 46810
rect 7733 46758 7779 46810
rect 7483 46756 7539 46758
rect 7563 46756 7619 46758
rect 7643 46756 7699 46758
rect 7723 46756 7779 46758
rect 7483 45722 7539 45724
rect 7563 45722 7619 45724
rect 7643 45722 7699 45724
rect 7723 45722 7779 45724
rect 7483 45670 7529 45722
rect 7529 45670 7539 45722
rect 7563 45670 7593 45722
rect 7593 45670 7605 45722
rect 7605 45670 7619 45722
rect 7643 45670 7657 45722
rect 7657 45670 7669 45722
rect 7669 45670 7699 45722
rect 7723 45670 7733 45722
rect 7733 45670 7779 45722
rect 7483 45668 7539 45670
rect 7563 45668 7619 45670
rect 7643 45668 7699 45670
rect 7723 45668 7779 45670
rect 7483 44634 7539 44636
rect 7563 44634 7619 44636
rect 7643 44634 7699 44636
rect 7723 44634 7779 44636
rect 7483 44582 7529 44634
rect 7529 44582 7539 44634
rect 7563 44582 7593 44634
rect 7593 44582 7605 44634
rect 7605 44582 7619 44634
rect 7643 44582 7657 44634
rect 7657 44582 7669 44634
rect 7669 44582 7699 44634
rect 7723 44582 7733 44634
rect 7733 44582 7779 44634
rect 7483 44580 7539 44582
rect 7563 44580 7619 44582
rect 7643 44580 7699 44582
rect 7723 44580 7779 44582
rect 7483 43546 7539 43548
rect 7563 43546 7619 43548
rect 7643 43546 7699 43548
rect 7723 43546 7779 43548
rect 7483 43494 7529 43546
rect 7529 43494 7539 43546
rect 7563 43494 7593 43546
rect 7593 43494 7605 43546
rect 7605 43494 7619 43546
rect 7643 43494 7657 43546
rect 7657 43494 7669 43546
rect 7669 43494 7699 43546
rect 7723 43494 7733 43546
rect 7733 43494 7779 43546
rect 7483 43492 7539 43494
rect 7563 43492 7619 43494
rect 7643 43492 7699 43494
rect 7723 43492 7779 43494
rect 7483 42458 7539 42460
rect 7563 42458 7619 42460
rect 7643 42458 7699 42460
rect 7723 42458 7779 42460
rect 7483 42406 7529 42458
rect 7529 42406 7539 42458
rect 7563 42406 7593 42458
rect 7593 42406 7605 42458
rect 7605 42406 7619 42458
rect 7643 42406 7657 42458
rect 7657 42406 7669 42458
rect 7669 42406 7699 42458
rect 7723 42406 7733 42458
rect 7733 42406 7779 42458
rect 7483 42404 7539 42406
rect 7563 42404 7619 42406
rect 7643 42404 7699 42406
rect 7723 42404 7779 42406
rect 7483 41370 7539 41372
rect 7563 41370 7619 41372
rect 7643 41370 7699 41372
rect 7723 41370 7779 41372
rect 7483 41318 7529 41370
rect 7529 41318 7539 41370
rect 7563 41318 7593 41370
rect 7593 41318 7605 41370
rect 7605 41318 7619 41370
rect 7643 41318 7657 41370
rect 7657 41318 7669 41370
rect 7669 41318 7699 41370
rect 7723 41318 7733 41370
rect 7733 41318 7779 41370
rect 7483 41316 7539 41318
rect 7563 41316 7619 41318
rect 7643 41316 7699 41318
rect 7723 41316 7779 41318
rect 7483 40282 7539 40284
rect 7563 40282 7619 40284
rect 7643 40282 7699 40284
rect 7723 40282 7779 40284
rect 7483 40230 7529 40282
rect 7529 40230 7539 40282
rect 7563 40230 7593 40282
rect 7593 40230 7605 40282
rect 7605 40230 7619 40282
rect 7643 40230 7657 40282
rect 7657 40230 7669 40282
rect 7669 40230 7699 40282
rect 7723 40230 7733 40282
rect 7733 40230 7779 40282
rect 7483 40228 7539 40230
rect 7563 40228 7619 40230
rect 7643 40228 7699 40230
rect 7723 40228 7779 40230
rect 7483 39194 7539 39196
rect 7563 39194 7619 39196
rect 7643 39194 7699 39196
rect 7723 39194 7779 39196
rect 7483 39142 7529 39194
rect 7529 39142 7539 39194
rect 7563 39142 7593 39194
rect 7593 39142 7605 39194
rect 7605 39142 7619 39194
rect 7643 39142 7657 39194
rect 7657 39142 7669 39194
rect 7669 39142 7699 39194
rect 7723 39142 7733 39194
rect 7733 39142 7779 39194
rect 7483 39140 7539 39142
rect 7563 39140 7619 39142
rect 7643 39140 7699 39142
rect 7723 39140 7779 39142
rect 7483 38106 7539 38108
rect 7563 38106 7619 38108
rect 7643 38106 7699 38108
rect 7723 38106 7779 38108
rect 7483 38054 7529 38106
rect 7529 38054 7539 38106
rect 7563 38054 7593 38106
rect 7593 38054 7605 38106
rect 7605 38054 7619 38106
rect 7643 38054 7657 38106
rect 7657 38054 7669 38106
rect 7669 38054 7699 38106
rect 7723 38054 7733 38106
rect 7733 38054 7779 38106
rect 7483 38052 7539 38054
rect 7563 38052 7619 38054
rect 7643 38052 7699 38054
rect 7723 38052 7779 38054
rect 7483 37018 7539 37020
rect 7563 37018 7619 37020
rect 7643 37018 7699 37020
rect 7723 37018 7779 37020
rect 7483 36966 7529 37018
rect 7529 36966 7539 37018
rect 7563 36966 7593 37018
rect 7593 36966 7605 37018
rect 7605 36966 7619 37018
rect 7643 36966 7657 37018
rect 7657 36966 7669 37018
rect 7669 36966 7699 37018
rect 7723 36966 7733 37018
rect 7733 36966 7779 37018
rect 7483 36964 7539 36966
rect 7563 36964 7619 36966
rect 7643 36964 7699 36966
rect 7723 36964 7779 36966
rect 7483 35930 7539 35932
rect 7563 35930 7619 35932
rect 7643 35930 7699 35932
rect 7723 35930 7779 35932
rect 7483 35878 7529 35930
rect 7529 35878 7539 35930
rect 7563 35878 7593 35930
rect 7593 35878 7605 35930
rect 7605 35878 7619 35930
rect 7643 35878 7657 35930
rect 7657 35878 7669 35930
rect 7669 35878 7699 35930
rect 7723 35878 7733 35930
rect 7733 35878 7779 35930
rect 7483 35876 7539 35878
rect 7563 35876 7619 35878
rect 7643 35876 7699 35878
rect 7723 35876 7779 35878
rect 7483 34842 7539 34844
rect 7563 34842 7619 34844
rect 7643 34842 7699 34844
rect 7723 34842 7779 34844
rect 7483 34790 7529 34842
rect 7529 34790 7539 34842
rect 7563 34790 7593 34842
rect 7593 34790 7605 34842
rect 7605 34790 7619 34842
rect 7643 34790 7657 34842
rect 7657 34790 7669 34842
rect 7669 34790 7699 34842
rect 7723 34790 7733 34842
rect 7733 34790 7779 34842
rect 7483 34788 7539 34790
rect 7563 34788 7619 34790
rect 7643 34788 7699 34790
rect 7723 34788 7779 34790
rect 7483 33754 7539 33756
rect 7563 33754 7619 33756
rect 7643 33754 7699 33756
rect 7723 33754 7779 33756
rect 7483 33702 7529 33754
rect 7529 33702 7539 33754
rect 7563 33702 7593 33754
rect 7593 33702 7605 33754
rect 7605 33702 7619 33754
rect 7643 33702 7657 33754
rect 7657 33702 7669 33754
rect 7669 33702 7699 33754
rect 7723 33702 7733 33754
rect 7733 33702 7779 33754
rect 7483 33700 7539 33702
rect 7563 33700 7619 33702
rect 7643 33700 7699 33702
rect 7723 33700 7779 33702
rect 7483 32666 7539 32668
rect 7563 32666 7619 32668
rect 7643 32666 7699 32668
rect 7723 32666 7779 32668
rect 7483 32614 7529 32666
rect 7529 32614 7539 32666
rect 7563 32614 7593 32666
rect 7593 32614 7605 32666
rect 7605 32614 7619 32666
rect 7643 32614 7657 32666
rect 7657 32614 7669 32666
rect 7669 32614 7699 32666
rect 7723 32614 7733 32666
rect 7733 32614 7779 32666
rect 7483 32612 7539 32614
rect 7563 32612 7619 32614
rect 7643 32612 7699 32614
rect 7723 32612 7779 32614
rect 7483 31578 7539 31580
rect 7563 31578 7619 31580
rect 7643 31578 7699 31580
rect 7723 31578 7779 31580
rect 7483 31526 7529 31578
rect 7529 31526 7539 31578
rect 7563 31526 7593 31578
rect 7593 31526 7605 31578
rect 7605 31526 7619 31578
rect 7643 31526 7657 31578
rect 7657 31526 7669 31578
rect 7669 31526 7699 31578
rect 7723 31526 7733 31578
rect 7733 31526 7779 31578
rect 7483 31524 7539 31526
rect 7563 31524 7619 31526
rect 7643 31524 7699 31526
rect 7723 31524 7779 31526
rect 7483 30490 7539 30492
rect 7563 30490 7619 30492
rect 7643 30490 7699 30492
rect 7723 30490 7779 30492
rect 7483 30438 7529 30490
rect 7529 30438 7539 30490
rect 7563 30438 7593 30490
rect 7593 30438 7605 30490
rect 7605 30438 7619 30490
rect 7643 30438 7657 30490
rect 7657 30438 7669 30490
rect 7669 30438 7699 30490
rect 7723 30438 7733 30490
rect 7733 30438 7779 30490
rect 7483 30436 7539 30438
rect 7563 30436 7619 30438
rect 7643 30436 7699 30438
rect 7723 30436 7779 30438
rect 7483 29402 7539 29404
rect 7563 29402 7619 29404
rect 7643 29402 7699 29404
rect 7723 29402 7779 29404
rect 7483 29350 7529 29402
rect 7529 29350 7539 29402
rect 7563 29350 7593 29402
rect 7593 29350 7605 29402
rect 7605 29350 7619 29402
rect 7643 29350 7657 29402
rect 7657 29350 7669 29402
rect 7669 29350 7699 29402
rect 7723 29350 7733 29402
rect 7733 29350 7779 29402
rect 7483 29348 7539 29350
rect 7563 29348 7619 29350
rect 7643 29348 7699 29350
rect 7723 29348 7779 29350
rect 7483 28314 7539 28316
rect 7563 28314 7619 28316
rect 7643 28314 7699 28316
rect 7723 28314 7779 28316
rect 7483 28262 7529 28314
rect 7529 28262 7539 28314
rect 7563 28262 7593 28314
rect 7593 28262 7605 28314
rect 7605 28262 7619 28314
rect 7643 28262 7657 28314
rect 7657 28262 7669 28314
rect 7669 28262 7699 28314
rect 7723 28262 7733 28314
rect 7733 28262 7779 28314
rect 7483 28260 7539 28262
rect 7563 28260 7619 28262
rect 7643 28260 7699 28262
rect 7723 28260 7779 28262
rect 7483 27226 7539 27228
rect 7563 27226 7619 27228
rect 7643 27226 7699 27228
rect 7723 27226 7779 27228
rect 7483 27174 7529 27226
rect 7529 27174 7539 27226
rect 7563 27174 7593 27226
rect 7593 27174 7605 27226
rect 7605 27174 7619 27226
rect 7643 27174 7657 27226
rect 7657 27174 7669 27226
rect 7669 27174 7699 27226
rect 7723 27174 7733 27226
rect 7733 27174 7779 27226
rect 7483 27172 7539 27174
rect 7563 27172 7619 27174
rect 7643 27172 7699 27174
rect 7723 27172 7779 27174
rect 7483 26138 7539 26140
rect 7563 26138 7619 26140
rect 7643 26138 7699 26140
rect 7723 26138 7779 26140
rect 7483 26086 7529 26138
rect 7529 26086 7539 26138
rect 7563 26086 7593 26138
rect 7593 26086 7605 26138
rect 7605 26086 7619 26138
rect 7643 26086 7657 26138
rect 7657 26086 7669 26138
rect 7669 26086 7699 26138
rect 7723 26086 7733 26138
rect 7733 26086 7779 26138
rect 7483 26084 7539 26086
rect 7563 26084 7619 26086
rect 7643 26084 7699 26086
rect 7723 26084 7779 26086
rect 7483 25050 7539 25052
rect 7563 25050 7619 25052
rect 7643 25050 7699 25052
rect 7723 25050 7779 25052
rect 7483 24998 7529 25050
rect 7529 24998 7539 25050
rect 7563 24998 7593 25050
rect 7593 24998 7605 25050
rect 7605 24998 7619 25050
rect 7643 24998 7657 25050
rect 7657 24998 7669 25050
rect 7669 24998 7699 25050
rect 7723 24998 7733 25050
rect 7733 24998 7779 25050
rect 7483 24996 7539 24998
rect 7563 24996 7619 24998
rect 7643 24996 7699 24998
rect 7723 24996 7779 24998
rect 7483 23962 7539 23964
rect 7563 23962 7619 23964
rect 7643 23962 7699 23964
rect 7723 23962 7779 23964
rect 7483 23910 7529 23962
rect 7529 23910 7539 23962
rect 7563 23910 7593 23962
rect 7593 23910 7605 23962
rect 7605 23910 7619 23962
rect 7643 23910 7657 23962
rect 7657 23910 7669 23962
rect 7669 23910 7699 23962
rect 7723 23910 7733 23962
rect 7733 23910 7779 23962
rect 7483 23908 7539 23910
rect 7563 23908 7619 23910
rect 7643 23908 7699 23910
rect 7723 23908 7779 23910
rect 7483 22874 7539 22876
rect 7563 22874 7619 22876
rect 7643 22874 7699 22876
rect 7723 22874 7779 22876
rect 7483 22822 7529 22874
rect 7529 22822 7539 22874
rect 7563 22822 7593 22874
rect 7593 22822 7605 22874
rect 7605 22822 7619 22874
rect 7643 22822 7657 22874
rect 7657 22822 7669 22874
rect 7669 22822 7699 22874
rect 7723 22822 7733 22874
rect 7733 22822 7779 22874
rect 7483 22820 7539 22822
rect 7563 22820 7619 22822
rect 7643 22820 7699 22822
rect 7723 22820 7779 22822
rect 7483 21786 7539 21788
rect 7563 21786 7619 21788
rect 7643 21786 7699 21788
rect 7723 21786 7779 21788
rect 7483 21734 7529 21786
rect 7529 21734 7539 21786
rect 7563 21734 7593 21786
rect 7593 21734 7605 21786
rect 7605 21734 7619 21786
rect 7643 21734 7657 21786
rect 7657 21734 7669 21786
rect 7669 21734 7699 21786
rect 7723 21734 7733 21786
rect 7733 21734 7779 21786
rect 7483 21732 7539 21734
rect 7563 21732 7619 21734
rect 7643 21732 7699 21734
rect 7723 21732 7779 21734
rect 7483 20698 7539 20700
rect 7563 20698 7619 20700
rect 7643 20698 7699 20700
rect 7723 20698 7779 20700
rect 7483 20646 7529 20698
rect 7529 20646 7539 20698
rect 7563 20646 7593 20698
rect 7593 20646 7605 20698
rect 7605 20646 7619 20698
rect 7643 20646 7657 20698
rect 7657 20646 7669 20698
rect 7669 20646 7699 20698
rect 7723 20646 7733 20698
rect 7733 20646 7779 20698
rect 7483 20644 7539 20646
rect 7563 20644 7619 20646
rect 7643 20644 7699 20646
rect 7723 20644 7779 20646
rect 7483 19610 7539 19612
rect 7563 19610 7619 19612
rect 7643 19610 7699 19612
rect 7723 19610 7779 19612
rect 7483 19558 7529 19610
rect 7529 19558 7539 19610
rect 7563 19558 7593 19610
rect 7593 19558 7605 19610
rect 7605 19558 7619 19610
rect 7643 19558 7657 19610
rect 7657 19558 7669 19610
rect 7669 19558 7699 19610
rect 7723 19558 7733 19610
rect 7733 19558 7779 19610
rect 7483 19556 7539 19558
rect 7563 19556 7619 19558
rect 7643 19556 7699 19558
rect 7723 19556 7779 19558
rect 7483 18522 7539 18524
rect 7563 18522 7619 18524
rect 7643 18522 7699 18524
rect 7723 18522 7779 18524
rect 7483 18470 7529 18522
rect 7529 18470 7539 18522
rect 7563 18470 7593 18522
rect 7593 18470 7605 18522
rect 7605 18470 7619 18522
rect 7643 18470 7657 18522
rect 7657 18470 7669 18522
rect 7669 18470 7699 18522
rect 7723 18470 7733 18522
rect 7733 18470 7779 18522
rect 7483 18468 7539 18470
rect 7563 18468 7619 18470
rect 7643 18468 7699 18470
rect 7723 18468 7779 18470
rect 7483 17434 7539 17436
rect 7563 17434 7619 17436
rect 7643 17434 7699 17436
rect 7723 17434 7779 17436
rect 7483 17382 7529 17434
rect 7529 17382 7539 17434
rect 7563 17382 7593 17434
rect 7593 17382 7605 17434
rect 7605 17382 7619 17434
rect 7643 17382 7657 17434
rect 7657 17382 7669 17434
rect 7669 17382 7699 17434
rect 7723 17382 7733 17434
rect 7733 17382 7779 17434
rect 7483 17380 7539 17382
rect 7563 17380 7619 17382
rect 7643 17380 7699 17382
rect 7723 17380 7779 17382
rect 7483 16346 7539 16348
rect 7563 16346 7619 16348
rect 7643 16346 7699 16348
rect 7723 16346 7779 16348
rect 7483 16294 7529 16346
rect 7529 16294 7539 16346
rect 7563 16294 7593 16346
rect 7593 16294 7605 16346
rect 7605 16294 7619 16346
rect 7643 16294 7657 16346
rect 7657 16294 7669 16346
rect 7669 16294 7699 16346
rect 7723 16294 7733 16346
rect 7733 16294 7779 16346
rect 7483 16292 7539 16294
rect 7563 16292 7619 16294
rect 7643 16292 7699 16294
rect 7723 16292 7779 16294
rect 7483 15258 7539 15260
rect 7563 15258 7619 15260
rect 7643 15258 7699 15260
rect 7723 15258 7779 15260
rect 7483 15206 7529 15258
rect 7529 15206 7539 15258
rect 7563 15206 7593 15258
rect 7593 15206 7605 15258
rect 7605 15206 7619 15258
rect 7643 15206 7657 15258
rect 7657 15206 7669 15258
rect 7669 15206 7699 15258
rect 7723 15206 7733 15258
rect 7733 15206 7779 15258
rect 7483 15204 7539 15206
rect 7563 15204 7619 15206
rect 7643 15204 7699 15206
rect 7723 15204 7779 15206
rect 7483 14170 7539 14172
rect 7563 14170 7619 14172
rect 7643 14170 7699 14172
rect 7723 14170 7779 14172
rect 7483 14118 7529 14170
rect 7529 14118 7539 14170
rect 7563 14118 7593 14170
rect 7593 14118 7605 14170
rect 7605 14118 7619 14170
rect 7643 14118 7657 14170
rect 7657 14118 7669 14170
rect 7669 14118 7699 14170
rect 7723 14118 7733 14170
rect 7733 14118 7779 14170
rect 7483 14116 7539 14118
rect 7563 14116 7619 14118
rect 7643 14116 7699 14118
rect 7723 14116 7779 14118
rect 7483 13082 7539 13084
rect 7563 13082 7619 13084
rect 7643 13082 7699 13084
rect 7723 13082 7779 13084
rect 7483 13030 7529 13082
rect 7529 13030 7539 13082
rect 7563 13030 7593 13082
rect 7593 13030 7605 13082
rect 7605 13030 7619 13082
rect 7643 13030 7657 13082
rect 7657 13030 7669 13082
rect 7669 13030 7699 13082
rect 7723 13030 7733 13082
rect 7733 13030 7779 13082
rect 7483 13028 7539 13030
rect 7563 13028 7619 13030
rect 7643 13028 7699 13030
rect 7723 13028 7779 13030
rect 7483 11994 7539 11996
rect 7563 11994 7619 11996
rect 7643 11994 7699 11996
rect 7723 11994 7779 11996
rect 7483 11942 7529 11994
rect 7529 11942 7539 11994
rect 7563 11942 7593 11994
rect 7593 11942 7605 11994
rect 7605 11942 7619 11994
rect 7643 11942 7657 11994
rect 7657 11942 7669 11994
rect 7669 11942 7699 11994
rect 7723 11942 7733 11994
rect 7733 11942 7779 11994
rect 7483 11940 7539 11942
rect 7563 11940 7619 11942
rect 7643 11940 7699 11942
rect 7723 11940 7779 11942
rect 7483 10906 7539 10908
rect 7563 10906 7619 10908
rect 7643 10906 7699 10908
rect 7723 10906 7779 10908
rect 7483 10854 7529 10906
rect 7529 10854 7539 10906
rect 7563 10854 7593 10906
rect 7593 10854 7605 10906
rect 7605 10854 7619 10906
rect 7643 10854 7657 10906
rect 7657 10854 7669 10906
rect 7669 10854 7699 10906
rect 7723 10854 7733 10906
rect 7733 10854 7779 10906
rect 7483 10852 7539 10854
rect 7563 10852 7619 10854
rect 7643 10852 7699 10854
rect 7723 10852 7779 10854
rect 7483 9818 7539 9820
rect 7563 9818 7619 9820
rect 7643 9818 7699 9820
rect 7723 9818 7779 9820
rect 7483 9766 7529 9818
rect 7529 9766 7539 9818
rect 7563 9766 7593 9818
rect 7593 9766 7605 9818
rect 7605 9766 7619 9818
rect 7643 9766 7657 9818
rect 7657 9766 7669 9818
rect 7669 9766 7699 9818
rect 7723 9766 7733 9818
rect 7733 9766 7779 9818
rect 7483 9764 7539 9766
rect 7563 9764 7619 9766
rect 7643 9764 7699 9766
rect 7723 9764 7779 9766
rect 7483 8730 7539 8732
rect 7563 8730 7619 8732
rect 7643 8730 7699 8732
rect 7723 8730 7779 8732
rect 7483 8678 7529 8730
rect 7529 8678 7539 8730
rect 7563 8678 7593 8730
rect 7593 8678 7605 8730
rect 7605 8678 7619 8730
rect 7643 8678 7657 8730
rect 7657 8678 7669 8730
rect 7669 8678 7699 8730
rect 7723 8678 7733 8730
rect 7733 8678 7779 8730
rect 7483 8676 7539 8678
rect 7563 8676 7619 8678
rect 7643 8676 7699 8678
rect 7723 8676 7779 8678
rect 5851 8186 5907 8188
rect 5931 8186 5987 8188
rect 6011 8186 6067 8188
rect 6091 8186 6147 8188
rect 5851 8134 5897 8186
rect 5897 8134 5907 8186
rect 5931 8134 5961 8186
rect 5961 8134 5973 8186
rect 5973 8134 5987 8186
rect 6011 8134 6025 8186
rect 6025 8134 6037 8186
rect 6037 8134 6067 8186
rect 6091 8134 6101 8186
rect 6101 8134 6147 8186
rect 5851 8132 5907 8134
rect 5931 8132 5987 8134
rect 6011 8132 6067 8134
rect 6091 8132 6147 8134
rect 7483 7642 7539 7644
rect 7563 7642 7619 7644
rect 7643 7642 7699 7644
rect 7723 7642 7779 7644
rect 7483 7590 7529 7642
rect 7529 7590 7539 7642
rect 7563 7590 7593 7642
rect 7593 7590 7605 7642
rect 7605 7590 7619 7642
rect 7643 7590 7657 7642
rect 7657 7590 7669 7642
rect 7669 7590 7699 7642
rect 7723 7590 7733 7642
rect 7733 7590 7779 7642
rect 7483 7588 7539 7590
rect 7563 7588 7619 7590
rect 7643 7588 7699 7590
rect 7723 7588 7779 7590
rect 5851 7098 5907 7100
rect 5931 7098 5987 7100
rect 6011 7098 6067 7100
rect 6091 7098 6147 7100
rect 5851 7046 5897 7098
rect 5897 7046 5907 7098
rect 5931 7046 5961 7098
rect 5961 7046 5973 7098
rect 5973 7046 5987 7098
rect 6011 7046 6025 7098
rect 6025 7046 6037 7098
rect 6037 7046 6067 7098
rect 6091 7046 6101 7098
rect 6101 7046 6147 7098
rect 5851 7044 5907 7046
rect 5931 7044 5987 7046
rect 6011 7044 6067 7046
rect 6091 7044 6147 7046
rect 10230 75656 10286 75712
rect 10138 74840 10194 74896
rect 9115 74554 9171 74556
rect 9195 74554 9251 74556
rect 9275 74554 9331 74556
rect 9355 74554 9411 74556
rect 9115 74502 9161 74554
rect 9161 74502 9171 74554
rect 9195 74502 9225 74554
rect 9225 74502 9237 74554
rect 9237 74502 9251 74554
rect 9275 74502 9289 74554
rect 9289 74502 9301 74554
rect 9301 74502 9331 74554
rect 9355 74502 9365 74554
rect 9365 74502 9411 74554
rect 9115 74500 9171 74502
rect 9195 74500 9251 74502
rect 9275 74500 9331 74502
rect 9355 74500 9411 74502
rect 9115 73466 9171 73468
rect 9195 73466 9251 73468
rect 9275 73466 9331 73468
rect 9355 73466 9411 73468
rect 9115 73414 9161 73466
rect 9161 73414 9171 73466
rect 9195 73414 9225 73466
rect 9225 73414 9237 73466
rect 9237 73414 9251 73466
rect 9275 73414 9289 73466
rect 9289 73414 9301 73466
rect 9301 73414 9331 73466
rect 9355 73414 9365 73466
rect 9365 73414 9411 73466
rect 9115 73412 9171 73414
rect 9195 73412 9251 73414
rect 9275 73412 9331 73414
rect 9355 73412 9411 73414
rect 9115 72378 9171 72380
rect 9195 72378 9251 72380
rect 9275 72378 9331 72380
rect 9355 72378 9411 72380
rect 9115 72326 9161 72378
rect 9161 72326 9171 72378
rect 9195 72326 9225 72378
rect 9225 72326 9237 72378
rect 9237 72326 9251 72378
rect 9275 72326 9289 72378
rect 9289 72326 9301 72378
rect 9301 72326 9331 72378
rect 9355 72326 9365 72378
rect 9365 72326 9411 72378
rect 9115 72324 9171 72326
rect 9195 72324 9251 72326
rect 9275 72324 9331 72326
rect 9355 72324 9411 72326
rect 10138 74024 10194 74080
rect 10138 73344 10194 73400
rect 10138 72528 10194 72584
rect 10138 71712 10194 71768
rect 9115 71290 9171 71292
rect 9195 71290 9251 71292
rect 9275 71290 9331 71292
rect 9355 71290 9411 71292
rect 9115 71238 9161 71290
rect 9161 71238 9171 71290
rect 9195 71238 9225 71290
rect 9225 71238 9237 71290
rect 9237 71238 9251 71290
rect 9275 71238 9289 71290
rect 9289 71238 9301 71290
rect 9301 71238 9331 71290
rect 9355 71238 9365 71290
rect 9365 71238 9411 71290
rect 9115 71236 9171 71238
rect 9195 71236 9251 71238
rect 9275 71236 9331 71238
rect 9355 71236 9411 71238
rect 10138 71032 10194 71088
rect 10138 70216 10194 70272
rect 9115 70202 9171 70204
rect 9195 70202 9251 70204
rect 9275 70202 9331 70204
rect 9355 70202 9411 70204
rect 9115 70150 9161 70202
rect 9161 70150 9171 70202
rect 9195 70150 9225 70202
rect 9225 70150 9237 70202
rect 9237 70150 9251 70202
rect 9275 70150 9289 70202
rect 9289 70150 9301 70202
rect 9301 70150 9331 70202
rect 9355 70150 9365 70202
rect 9365 70150 9411 70202
rect 9115 70148 9171 70150
rect 9195 70148 9251 70150
rect 9275 70148 9331 70150
rect 9355 70148 9411 70150
rect 10138 69400 10194 69456
rect 9115 69114 9171 69116
rect 9195 69114 9251 69116
rect 9275 69114 9331 69116
rect 9355 69114 9411 69116
rect 9115 69062 9161 69114
rect 9161 69062 9171 69114
rect 9195 69062 9225 69114
rect 9225 69062 9237 69114
rect 9237 69062 9251 69114
rect 9275 69062 9289 69114
rect 9289 69062 9301 69114
rect 9301 69062 9331 69114
rect 9355 69062 9365 69114
rect 9365 69062 9411 69114
rect 9115 69060 9171 69062
rect 9195 69060 9251 69062
rect 9275 69060 9331 69062
rect 9355 69060 9411 69062
rect 10138 68756 10140 68776
rect 10140 68756 10192 68776
rect 10192 68756 10194 68776
rect 10138 68720 10194 68756
rect 9115 68026 9171 68028
rect 9195 68026 9251 68028
rect 9275 68026 9331 68028
rect 9355 68026 9411 68028
rect 9115 67974 9161 68026
rect 9161 67974 9171 68026
rect 9195 67974 9225 68026
rect 9225 67974 9237 68026
rect 9237 67974 9251 68026
rect 9275 67974 9289 68026
rect 9289 67974 9301 68026
rect 9301 67974 9331 68026
rect 9355 67974 9365 68026
rect 9365 67974 9411 68026
rect 9115 67972 9171 67974
rect 9195 67972 9251 67974
rect 9275 67972 9331 67974
rect 9355 67972 9411 67974
rect 10138 67904 10194 67960
rect 10138 67088 10194 67144
rect 9115 66938 9171 66940
rect 9195 66938 9251 66940
rect 9275 66938 9331 66940
rect 9355 66938 9411 66940
rect 9115 66886 9161 66938
rect 9161 66886 9171 66938
rect 9195 66886 9225 66938
rect 9225 66886 9237 66938
rect 9237 66886 9251 66938
rect 9275 66886 9289 66938
rect 9289 66886 9301 66938
rect 9301 66886 9331 66938
rect 9355 66886 9365 66938
rect 9365 66886 9411 66938
rect 9115 66884 9171 66886
rect 9195 66884 9251 66886
rect 9275 66884 9331 66886
rect 9355 66884 9411 66886
rect 9115 65850 9171 65852
rect 9195 65850 9251 65852
rect 9275 65850 9331 65852
rect 9355 65850 9411 65852
rect 9115 65798 9161 65850
rect 9161 65798 9171 65850
rect 9195 65798 9225 65850
rect 9225 65798 9237 65850
rect 9237 65798 9251 65850
rect 9275 65798 9289 65850
rect 9289 65798 9301 65850
rect 9301 65798 9331 65850
rect 9355 65798 9365 65850
rect 9365 65798 9411 65850
rect 9115 65796 9171 65798
rect 9195 65796 9251 65798
rect 9275 65796 9331 65798
rect 9355 65796 9411 65798
rect 10138 66408 10194 66464
rect 10138 65592 10194 65648
rect 10138 64776 10194 64832
rect 9115 64762 9171 64764
rect 9195 64762 9251 64764
rect 9275 64762 9331 64764
rect 9355 64762 9411 64764
rect 9115 64710 9161 64762
rect 9161 64710 9171 64762
rect 9195 64710 9225 64762
rect 9225 64710 9237 64762
rect 9237 64710 9251 64762
rect 9275 64710 9289 64762
rect 9289 64710 9301 64762
rect 9301 64710 9331 64762
rect 9355 64710 9365 64762
rect 9365 64710 9411 64762
rect 9115 64708 9171 64710
rect 9195 64708 9251 64710
rect 9275 64708 9331 64710
rect 9355 64708 9411 64710
rect 9115 63674 9171 63676
rect 9195 63674 9251 63676
rect 9275 63674 9331 63676
rect 9355 63674 9411 63676
rect 9115 63622 9161 63674
rect 9161 63622 9171 63674
rect 9195 63622 9225 63674
rect 9225 63622 9237 63674
rect 9237 63622 9251 63674
rect 9275 63622 9289 63674
rect 9289 63622 9301 63674
rect 9301 63622 9331 63674
rect 9355 63622 9365 63674
rect 9365 63622 9411 63674
rect 9115 63620 9171 63622
rect 9195 63620 9251 63622
rect 9275 63620 9331 63622
rect 9355 63620 9411 63622
rect 9115 62586 9171 62588
rect 9195 62586 9251 62588
rect 9275 62586 9331 62588
rect 9355 62586 9411 62588
rect 9115 62534 9161 62586
rect 9161 62534 9171 62586
rect 9195 62534 9225 62586
rect 9225 62534 9237 62586
rect 9237 62534 9251 62586
rect 9275 62534 9289 62586
rect 9289 62534 9301 62586
rect 9301 62534 9331 62586
rect 9355 62534 9365 62586
rect 9365 62534 9411 62586
rect 9115 62532 9171 62534
rect 9195 62532 9251 62534
rect 9275 62532 9331 62534
rect 9355 62532 9411 62534
rect 9115 61498 9171 61500
rect 9195 61498 9251 61500
rect 9275 61498 9331 61500
rect 9355 61498 9411 61500
rect 9115 61446 9161 61498
rect 9161 61446 9171 61498
rect 9195 61446 9225 61498
rect 9225 61446 9237 61498
rect 9237 61446 9251 61498
rect 9275 61446 9289 61498
rect 9289 61446 9301 61498
rect 9301 61446 9331 61498
rect 9355 61446 9365 61498
rect 9365 61446 9411 61498
rect 9115 61444 9171 61446
rect 9195 61444 9251 61446
rect 9275 61444 9331 61446
rect 9355 61444 9411 61446
rect 9115 60410 9171 60412
rect 9195 60410 9251 60412
rect 9275 60410 9331 60412
rect 9355 60410 9411 60412
rect 9115 60358 9161 60410
rect 9161 60358 9171 60410
rect 9195 60358 9225 60410
rect 9225 60358 9237 60410
rect 9237 60358 9251 60410
rect 9275 60358 9289 60410
rect 9289 60358 9301 60410
rect 9301 60358 9331 60410
rect 9355 60358 9365 60410
rect 9365 60358 9411 60410
rect 9115 60356 9171 60358
rect 9195 60356 9251 60358
rect 9275 60356 9331 60358
rect 9355 60356 9411 60358
rect 10138 64096 10194 64152
rect 10138 63316 10140 63336
rect 10140 63316 10192 63336
rect 10192 63316 10194 63336
rect 10138 63280 10194 63316
rect 10138 62464 10194 62520
rect 10138 61784 10194 61840
rect 10138 60968 10194 61024
rect 9115 59322 9171 59324
rect 9195 59322 9251 59324
rect 9275 59322 9331 59324
rect 9355 59322 9411 59324
rect 9115 59270 9161 59322
rect 9161 59270 9171 59322
rect 9195 59270 9225 59322
rect 9225 59270 9237 59322
rect 9237 59270 9251 59322
rect 9275 59270 9289 59322
rect 9289 59270 9301 59322
rect 9301 59270 9331 59322
rect 9355 59270 9365 59322
rect 9365 59270 9411 59322
rect 9115 59268 9171 59270
rect 9195 59268 9251 59270
rect 9275 59268 9331 59270
rect 9355 59268 9411 59270
rect 10138 60288 10194 60344
rect 10138 59472 10194 59528
rect 9115 58234 9171 58236
rect 9195 58234 9251 58236
rect 9275 58234 9331 58236
rect 9355 58234 9411 58236
rect 9115 58182 9161 58234
rect 9161 58182 9171 58234
rect 9195 58182 9225 58234
rect 9225 58182 9237 58234
rect 9237 58182 9251 58234
rect 9275 58182 9289 58234
rect 9289 58182 9301 58234
rect 9301 58182 9331 58234
rect 9355 58182 9365 58234
rect 9365 58182 9411 58234
rect 9115 58180 9171 58182
rect 9195 58180 9251 58182
rect 9275 58180 9331 58182
rect 9355 58180 9411 58182
rect 10138 58656 10194 58712
rect 10138 57976 10194 58032
rect 10138 57160 10194 57216
rect 9115 57146 9171 57148
rect 9195 57146 9251 57148
rect 9275 57146 9331 57148
rect 9355 57146 9411 57148
rect 9115 57094 9161 57146
rect 9161 57094 9171 57146
rect 9195 57094 9225 57146
rect 9225 57094 9237 57146
rect 9237 57094 9251 57146
rect 9275 57094 9289 57146
rect 9289 57094 9301 57146
rect 9301 57094 9331 57146
rect 9355 57094 9365 57146
rect 9365 57094 9411 57146
rect 9115 57092 9171 57094
rect 9195 57092 9251 57094
rect 9275 57092 9331 57094
rect 9355 57092 9411 57094
rect 10138 56344 10194 56400
rect 9115 56058 9171 56060
rect 9195 56058 9251 56060
rect 9275 56058 9331 56060
rect 9355 56058 9411 56060
rect 9115 56006 9161 56058
rect 9161 56006 9171 56058
rect 9195 56006 9225 56058
rect 9225 56006 9237 56058
rect 9237 56006 9251 56058
rect 9275 56006 9289 56058
rect 9289 56006 9301 56058
rect 9301 56006 9331 56058
rect 9355 56006 9365 56058
rect 9365 56006 9411 56058
rect 9115 56004 9171 56006
rect 9195 56004 9251 56006
rect 9275 56004 9331 56006
rect 9355 56004 9411 56006
rect 9115 54970 9171 54972
rect 9195 54970 9251 54972
rect 9275 54970 9331 54972
rect 9355 54970 9411 54972
rect 9115 54918 9161 54970
rect 9161 54918 9171 54970
rect 9195 54918 9225 54970
rect 9225 54918 9237 54970
rect 9237 54918 9251 54970
rect 9275 54918 9289 54970
rect 9289 54918 9301 54970
rect 9301 54918 9331 54970
rect 9355 54918 9365 54970
rect 9365 54918 9411 54970
rect 9115 54916 9171 54918
rect 9195 54916 9251 54918
rect 9275 54916 9331 54918
rect 9355 54916 9411 54918
rect 10138 55700 10140 55720
rect 10140 55700 10192 55720
rect 10192 55700 10194 55720
rect 10138 55664 10194 55700
rect 9115 53882 9171 53884
rect 9195 53882 9251 53884
rect 9275 53882 9331 53884
rect 9355 53882 9411 53884
rect 9115 53830 9161 53882
rect 9161 53830 9171 53882
rect 9195 53830 9225 53882
rect 9225 53830 9237 53882
rect 9237 53830 9251 53882
rect 9275 53830 9289 53882
rect 9289 53830 9301 53882
rect 9301 53830 9331 53882
rect 9355 53830 9365 53882
rect 9365 53830 9411 53882
rect 9115 53828 9171 53830
rect 9195 53828 9251 53830
rect 9275 53828 9331 53830
rect 9355 53828 9411 53830
rect 10230 54848 10286 54904
rect 10046 54052 10102 54088
rect 10046 54032 10048 54052
rect 10048 54032 10100 54052
rect 10100 54032 10102 54052
rect 10046 53388 10048 53408
rect 10048 53388 10100 53408
rect 10100 53388 10102 53408
rect 10046 53352 10102 53388
rect 9115 52794 9171 52796
rect 9195 52794 9251 52796
rect 9275 52794 9331 52796
rect 9355 52794 9411 52796
rect 9115 52742 9161 52794
rect 9161 52742 9171 52794
rect 9195 52742 9225 52794
rect 9225 52742 9237 52794
rect 9237 52742 9251 52794
rect 9275 52742 9289 52794
rect 9289 52742 9301 52794
rect 9301 52742 9331 52794
rect 9355 52742 9365 52794
rect 9365 52742 9411 52794
rect 9115 52740 9171 52742
rect 9195 52740 9251 52742
rect 9275 52740 9331 52742
rect 9355 52740 9411 52742
rect 10046 52536 10102 52592
rect 10046 51756 10048 51776
rect 10048 51756 10100 51776
rect 10100 51756 10102 51776
rect 10046 51720 10102 51756
rect 9115 51706 9171 51708
rect 9195 51706 9251 51708
rect 9275 51706 9331 51708
rect 9355 51706 9411 51708
rect 9115 51654 9161 51706
rect 9161 51654 9171 51706
rect 9195 51654 9225 51706
rect 9225 51654 9237 51706
rect 9237 51654 9251 51706
rect 9275 51654 9289 51706
rect 9289 51654 9301 51706
rect 9301 51654 9331 51706
rect 9355 51654 9365 51706
rect 9365 51654 9411 51706
rect 9115 51652 9171 51654
rect 9195 51652 9251 51654
rect 9275 51652 9331 51654
rect 9355 51652 9411 51654
rect 10046 51040 10102 51096
rect 9115 50618 9171 50620
rect 9195 50618 9251 50620
rect 9275 50618 9331 50620
rect 9355 50618 9411 50620
rect 9115 50566 9161 50618
rect 9161 50566 9171 50618
rect 9195 50566 9225 50618
rect 9225 50566 9237 50618
rect 9237 50566 9251 50618
rect 9275 50566 9289 50618
rect 9289 50566 9301 50618
rect 9301 50566 9331 50618
rect 9355 50566 9365 50618
rect 9365 50566 9411 50618
rect 9115 50564 9171 50566
rect 9195 50564 9251 50566
rect 9275 50564 9331 50566
rect 9355 50564 9411 50566
rect 10046 50224 10102 50280
rect 9115 49530 9171 49532
rect 9195 49530 9251 49532
rect 9275 49530 9331 49532
rect 9355 49530 9411 49532
rect 9115 49478 9161 49530
rect 9161 49478 9171 49530
rect 9195 49478 9225 49530
rect 9225 49478 9237 49530
rect 9237 49478 9251 49530
rect 9275 49478 9289 49530
rect 9289 49478 9301 49530
rect 9301 49478 9331 49530
rect 9355 49478 9365 49530
rect 9365 49478 9411 49530
rect 9115 49476 9171 49478
rect 9195 49476 9251 49478
rect 9275 49476 9331 49478
rect 9355 49476 9411 49478
rect 9115 48442 9171 48444
rect 9195 48442 9251 48444
rect 9275 48442 9331 48444
rect 9355 48442 9411 48444
rect 9115 48390 9161 48442
rect 9161 48390 9171 48442
rect 9195 48390 9225 48442
rect 9225 48390 9237 48442
rect 9237 48390 9251 48442
rect 9275 48390 9289 48442
rect 9289 48390 9301 48442
rect 9301 48390 9331 48442
rect 9355 48390 9365 48442
rect 9365 48390 9411 48442
rect 9115 48388 9171 48390
rect 9195 48388 9251 48390
rect 9275 48388 9331 48390
rect 9355 48388 9411 48390
rect 9115 47354 9171 47356
rect 9195 47354 9251 47356
rect 9275 47354 9331 47356
rect 9355 47354 9411 47356
rect 9115 47302 9161 47354
rect 9161 47302 9171 47354
rect 9195 47302 9225 47354
rect 9225 47302 9237 47354
rect 9237 47302 9251 47354
rect 9275 47302 9289 47354
rect 9289 47302 9301 47354
rect 9301 47302 9331 47354
rect 9355 47302 9365 47354
rect 9365 47302 9411 47354
rect 9115 47300 9171 47302
rect 9195 47300 9251 47302
rect 9275 47300 9331 47302
rect 9355 47300 9411 47302
rect 10046 49408 10102 49464
rect 10046 48728 10102 48784
rect 10046 47948 10048 47968
rect 10048 47948 10100 47968
rect 10100 47948 10102 47968
rect 10046 47912 10102 47948
rect 10046 47096 10102 47152
rect 10046 46436 10102 46472
rect 10046 46416 10048 46436
rect 10048 46416 10100 46436
rect 10100 46416 10102 46436
rect 9115 46266 9171 46268
rect 9195 46266 9251 46268
rect 9275 46266 9331 46268
rect 9355 46266 9411 46268
rect 9115 46214 9161 46266
rect 9161 46214 9171 46266
rect 9195 46214 9225 46266
rect 9225 46214 9237 46266
rect 9237 46214 9251 46266
rect 9275 46214 9289 46266
rect 9289 46214 9301 46266
rect 9301 46214 9331 46266
rect 9355 46214 9365 46266
rect 9365 46214 9411 46266
rect 9115 46212 9171 46214
rect 9195 46212 9251 46214
rect 9275 46212 9331 46214
rect 9355 46212 9411 46214
rect 9115 45178 9171 45180
rect 9195 45178 9251 45180
rect 9275 45178 9331 45180
rect 9355 45178 9411 45180
rect 9115 45126 9161 45178
rect 9161 45126 9171 45178
rect 9195 45126 9225 45178
rect 9225 45126 9237 45178
rect 9237 45126 9251 45178
rect 9275 45126 9289 45178
rect 9289 45126 9301 45178
rect 9301 45126 9331 45178
rect 9355 45126 9365 45178
rect 9365 45126 9411 45178
rect 9115 45124 9171 45126
rect 9195 45124 9251 45126
rect 9275 45124 9331 45126
rect 9355 45124 9411 45126
rect 9115 44090 9171 44092
rect 9195 44090 9251 44092
rect 9275 44090 9331 44092
rect 9355 44090 9411 44092
rect 9115 44038 9161 44090
rect 9161 44038 9171 44090
rect 9195 44038 9225 44090
rect 9225 44038 9237 44090
rect 9237 44038 9251 44090
rect 9275 44038 9289 44090
rect 9289 44038 9301 44090
rect 9301 44038 9331 44090
rect 9355 44038 9365 44090
rect 9365 44038 9411 44090
rect 9115 44036 9171 44038
rect 9195 44036 9251 44038
rect 9275 44036 9331 44038
rect 9355 44036 9411 44038
rect 9115 43002 9171 43004
rect 9195 43002 9251 43004
rect 9275 43002 9331 43004
rect 9355 43002 9411 43004
rect 9115 42950 9161 43002
rect 9161 42950 9171 43002
rect 9195 42950 9225 43002
rect 9225 42950 9237 43002
rect 9237 42950 9251 43002
rect 9275 42950 9289 43002
rect 9289 42950 9301 43002
rect 9301 42950 9331 43002
rect 9355 42950 9365 43002
rect 9365 42950 9411 43002
rect 9115 42948 9171 42950
rect 9195 42948 9251 42950
rect 9275 42948 9331 42950
rect 9355 42948 9411 42950
rect 10046 45600 10102 45656
rect 10046 44784 10102 44840
rect 10046 44140 10048 44160
rect 10048 44140 10100 44160
rect 10100 44140 10102 44160
rect 10046 44104 10102 44140
rect 10046 43288 10102 43344
rect 10046 42508 10048 42528
rect 10048 42508 10100 42528
rect 10100 42508 10102 42528
rect 10046 42472 10102 42508
rect 9115 41914 9171 41916
rect 9195 41914 9251 41916
rect 9275 41914 9331 41916
rect 9355 41914 9411 41916
rect 9115 41862 9161 41914
rect 9161 41862 9171 41914
rect 9195 41862 9225 41914
rect 9225 41862 9237 41914
rect 9237 41862 9251 41914
rect 9275 41862 9289 41914
rect 9289 41862 9301 41914
rect 9301 41862 9331 41914
rect 9355 41862 9365 41914
rect 9365 41862 9411 41914
rect 9115 41860 9171 41862
rect 9195 41860 9251 41862
rect 9275 41860 9331 41862
rect 9355 41860 9411 41862
rect 10046 41792 10102 41848
rect 9115 40826 9171 40828
rect 9195 40826 9251 40828
rect 9275 40826 9331 40828
rect 9355 40826 9411 40828
rect 9115 40774 9161 40826
rect 9161 40774 9171 40826
rect 9195 40774 9225 40826
rect 9225 40774 9237 40826
rect 9237 40774 9251 40826
rect 9275 40774 9289 40826
rect 9289 40774 9301 40826
rect 9301 40774 9331 40826
rect 9355 40774 9365 40826
rect 9365 40774 9411 40826
rect 9115 40772 9171 40774
rect 9195 40772 9251 40774
rect 9275 40772 9331 40774
rect 9355 40772 9411 40774
rect 10046 40996 10102 41032
rect 10046 40976 10048 40996
rect 10048 40976 10100 40996
rect 10100 40976 10102 40996
rect 9115 39738 9171 39740
rect 9195 39738 9251 39740
rect 9275 39738 9331 39740
rect 9355 39738 9411 39740
rect 9115 39686 9161 39738
rect 9161 39686 9171 39738
rect 9195 39686 9225 39738
rect 9225 39686 9237 39738
rect 9237 39686 9251 39738
rect 9275 39686 9289 39738
rect 9289 39686 9301 39738
rect 9301 39686 9331 39738
rect 9355 39686 9365 39738
rect 9365 39686 9411 39738
rect 9115 39684 9171 39686
rect 9195 39684 9251 39686
rect 9275 39684 9331 39686
rect 9355 39684 9411 39686
rect 9115 38650 9171 38652
rect 9195 38650 9251 38652
rect 9275 38650 9331 38652
rect 9355 38650 9411 38652
rect 9115 38598 9161 38650
rect 9161 38598 9171 38650
rect 9195 38598 9225 38650
rect 9225 38598 9237 38650
rect 9237 38598 9251 38650
rect 9275 38598 9289 38650
rect 9289 38598 9301 38650
rect 9301 38598 9331 38650
rect 9355 38598 9365 38650
rect 9365 38598 9411 38650
rect 9115 38596 9171 38598
rect 9195 38596 9251 38598
rect 9275 38596 9331 38598
rect 9355 38596 9411 38598
rect 10046 40332 10048 40352
rect 10048 40332 10100 40352
rect 10100 40332 10102 40352
rect 10046 40296 10102 40332
rect 10046 39480 10102 39536
rect 9115 37562 9171 37564
rect 9195 37562 9251 37564
rect 9275 37562 9331 37564
rect 9355 37562 9411 37564
rect 9115 37510 9161 37562
rect 9161 37510 9171 37562
rect 9195 37510 9225 37562
rect 9225 37510 9237 37562
rect 9237 37510 9251 37562
rect 9275 37510 9289 37562
rect 9289 37510 9301 37562
rect 9301 37510 9331 37562
rect 9355 37510 9365 37562
rect 9365 37510 9411 37562
rect 9115 37508 9171 37510
rect 9195 37508 9251 37510
rect 9275 37508 9331 37510
rect 9355 37508 9411 37510
rect 10046 38700 10048 38720
rect 10048 38700 10100 38720
rect 10100 38700 10102 38720
rect 10046 38664 10102 38700
rect 10046 37984 10102 38040
rect 10046 37168 10102 37224
rect 9115 36474 9171 36476
rect 9195 36474 9251 36476
rect 9275 36474 9331 36476
rect 9355 36474 9411 36476
rect 9115 36422 9161 36474
rect 9161 36422 9171 36474
rect 9195 36422 9225 36474
rect 9225 36422 9237 36474
rect 9237 36422 9251 36474
rect 9275 36422 9289 36474
rect 9289 36422 9301 36474
rect 9301 36422 9331 36474
rect 9355 36422 9365 36474
rect 9365 36422 9411 36474
rect 9115 36420 9171 36422
rect 9195 36420 9251 36422
rect 9275 36420 9331 36422
rect 9355 36420 9411 36422
rect 9115 35386 9171 35388
rect 9195 35386 9251 35388
rect 9275 35386 9331 35388
rect 9355 35386 9411 35388
rect 9115 35334 9161 35386
rect 9161 35334 9171 35386
rect 9195 35334 9225 35386
rect 9225 35334 9237 35386
rect 9237 35334 9251 35386
rect 9275 35334 9289 35386
rect 9289 35334 9301 35386
rect 9301 35334 9331 35386
rect 9355 35334 9365 35386
rect 9365 35334 9411 35386
rect 9115 35332 9171 35334
rect 9195 35332 9251 35334
rect 9275 35332 9331 35334
rect 9355 35332 9411 35334
rect 9115 34298 9171 34300
rect 9195 34298 9251 34300
rect 9275 34298 9331 34300
rect 9355 34298 9411 34300
rect 9115 34246 9161 34298
rect 9161 34246 9171 34298
rect 9195 34246 9225 34298
rect 9225 34246 9237 34298
rect 9237 34246 9251 34298
rect 9275 34246 9289 34298
rect 9289 34246 9301 34298
rect 9301 34246 9331 34298
rect 9355 34246 9365 34298
rect 9365 34246 9411 34298
rect 9115 34244 9171 34246
rect 9195 34244 9251 34246
rect 9275 34244 9331 34246
rect 9355 34244 9411 34246
rect 9115 33210 9171 33212
rect 9195 33210 9251 33212
rect 9275 33210 9331 33212
rect 9355 33210 9411 33212
rect 9115 33158 9161 33210
rect 9161 33158 9171 33210
rect 9195 33158 9225 33210
rect 9225 33158 9237 33210
rect 9237 33158 9251 33210
rect 9275 33158 9289 33210
rect 9289 33158 9301 33210
rect 9301 33158 9331 33210
rect 9355 33158 9365 33210
rect 9365 33158 9411 33210
rect 9115 33156 9171 33158
rect 9195 33156 9251 33158
rect 9275 33156 9331 33158
rect 9355 33156 9411 33158
rect 10046 36352 10102 36408
rect 10046 35672 10102 35728
rect 10046 34892 10048 34912
rect 10048 34892 10100 34912
rect 10100 34892 10102 34912
rect 10046 34856 10102 34892
rect 10046 34040 10102 34096
rect 10046 33380 10102 33416
rect 10046 33360 10048 33380
rect 10048 33360 10100 33380
rect 10100 33360 10102 33380
rect 10046 32544 10102 32600
rect 9115 32122 9171 32124
rect 9195 32122 9251 32124
rect 9275 32122 9331 32124
rect 9355 32122 9411 32124
rect 9115 32070 9161 32122
rect 9161 32070 9171 32122
rect 9195 32070 9225 32122
rect 9225 32070 9237 32122
rect 9237 32070 9251 32122
rect 9275 32070 9289 32122
rect 9289 32070 9301 32122
rect 9301 32070 9331 32122
rect 9355 32070 9365 32122
rect 9365 32070 9411 32122
rect 9115 32068 9171 32070
rect 9195 32068 9251 32070
rect 9275 32068 9331 32070
rect 9355 32068 9411 32070
rect 10046 31728 10102 31784
rect 10046 31084 10048 31104
rect 10048 31084 10100 31104
rect 10100 31084 10102 31104
rect 10046 31048 10102 31084
rect 9115 31034 9171 31036
rect 9195 31034 9251 31036
rect 9275 31034 9331 31036
rect 9355 31034 9411 31036
rect 9115 30982 9161 31034
rect 9161 30982 9171 31034
rect 9195 30982 9225 31034
rect 9225 30982 9237 31034
rect 9237 30982 9251 31034
rect 9275 30982 9289 31034
rect 9289 30982 9301 31034
rect 9301 30982 9331 31034
rect 9355 30982 9365 31034
rect 9365 30982 9411 31034
rect 9115 30980 9171 30982
rect 9195 30980 9251 30982
rect 9275 30980 9331 30982
rect 9355 30980 9411 30982
rect 9115 29946 9171 29948
rect 9195 29946 9251 29948
rect 9275 29946 9331 29948
rect 9355 29946 9411 29948
rect 9115 29894 9161 29946
rect 9161 29894 9171 29946
rect 9195 29894 9225 29946
rect 9225 29894 9237 29946
rect 9237 29894 9251 29946
rect 9275 29894 9289 29946
rect 9289 29894 9301 29946
rect 9301 29894 9331 29946
rect 9355 29894 9365 29946
rect 9365 29894 9411 29946
rect 9115 29892 9171 29894
rect 9195 29892 9251 29894
rect 9275 29892 9331 29894
rect 9355 29892 9411 29894
rect 10046 30232 10102 30288
rect 9494 29416 9550 29472
rect 9115 28858 9171 28860
rect 9195 28858 9251 28860
rect 9275 28858 9331 28860
rect 9355 28858 9411 28860
rect 9115 28806 9161 28858
rect 9161 28806 9171 28858
rect 9195 28806 9225 28858
rect 9225 28806 9237 28858
rect 9237 28806 9251 28858
rect 9275 28806 9289 28858
rect 9289 28806 9301 28858
rect 9301 28806 9331 28858
rect 9355 28806 9365 28858
rect 9365 28806 9411 28858
rect 9115 28804 9171 28806
rect 9195 28804 9251 28806
rect 9275 28804 9331 28806
rect 9355 28804 9411 28806
rect 10138 28736 10194 28792
rect 10138 27920 10194 27976
rect 9115 27770 9171 27772
rect 9195 27770 9251 27772
rect 9275 27770 9331 27772
rect 9355 27770 9411 27772
rect 9115 27718 9161 27770
rect 9161 27718 9171 27770
rect 9195 27718 9225 27770
rect 9225 27718 9237 27770
rect 9237 27718 9251 27770
rect 9275 27718 9289 27770
rect 9289 27718 9301 27770
rect 9301 27718 9331 27770
rect 9355 27718 9365 27770
rect 9365 27718 9411 27770
rect 9115 27716 9171 27718
rect 9195 27716 9251 27718
rect 9275 27716 9331 27718
rect 9355 27716 9411 27718
rect 10138 27104 10194 27160
rect 9115 26682 9171 26684
rect 9195 26682 9251 26684
rect 9275 26682 9331 26684
rect 9355 26682 9411 26684
rect 9115 26630 9161 26682
rect 9161 26630 9171 26682
rect 9195 26630 9225 26682
rect 9225 26630 9237 26682
rect 9237 26630 9251 26682
rect 9275 26630 9289 26682
rect 9289 26630 9301 26682
rect 9301 26630 9331 26682
rect 9355 26630 9365 26682
rect 9365 26630 9411 26682
rect 9115 26628 9171 26630
rect 9195 26628 9251 26630
rect 9275 26628 9331 26630
rect 9355 26628 9411 26630
rect 10138 26444 10194 26480
rect 10138 26424 10140 26444
rect 10140 26424 10192 26444
rect 10192 26424 10194 26444
rect 10138 25608 10194 25664
rect 9115 25594 9171 25596
rect 9195 25594 9251 25596
rect 9275 25594 9331 25596
rect 9355 25594 9411 25596
rect 9115 25542 9161 25594
rect 9161 25542 9171 25594
rect 9195 25542 9225 25594
rect 9225 25542 9237 25594
rect 9237 25542 9251 25594
rect 9275 25542 9289 25594
rect 9289 25542 9301 25594
rect 9301 25542 9331 25594
rect 9355 25542 9365 25594
rect 9365 25542 9411 25594
rect 9115 25540 9171 25542
rect 9195 25540 9251 25542
rect 9275 25540 9331 25542
rect 9355 25540 9411 25542
rect 10138 24812 10194 24848
rect 10138 24792 10140 24812
rect 10140 24792 10192 24812
rect 10192 24792 10194 24812
rect 9115 24506 9171 24508
rect 9195 24506 9251 24508
rect 9275 24506 9331 24508
rect 9355 24506 9411 24508
rect 9115 24454 9161 24506
rect 9161 24454 9171 24506
rect 9195 24454 9225 24506
rect 9225 24454 9237 24506
rect 9237 24454 9251 24506
rect 9275 24454 9289 24506
rect 9289 24454 9301 24506
rect 9301 24454 9331 24506
rect 9355 24454 9365 24506
rect 9365 24454 9411 24506
rect 9115 24452 9171 24454
rect 9195 24452 9251 24454
rect 9275 24452 9331 24454
rect 9355 24452 9411 24454
rect 10138 24112 10194 24168
rect 9115 23418 9171 23420
rect 9195 23418 9251 23420
rect 9275 23418 9331 23420
rect 9355 23418 9411 23420
rect 9115 23366 9161 23418
rect 9161 23366 9171 23418
rect 9195 23366 9225 23418
rect 9225 23366 9237 23418
rect 9237 23366 9251 23418
rect 9275 23366 9289 23418
rect 9289 23366 9301 23418
rect 9301 23366 9331 23418
rect 9355 23366 9365 23418
rect 9365 23366 9411 23418
rect 9115 23364 9171 23366
rect 9195 23364 9251 23366
rect 9275 23364 9331 23366
rect 9355 23364 9411 23366
rect 10046 23296 10102 23352
rect 9115 22330 9171 22332
rect 9195 22330 9251 22332
rect 9275 22330 9331 22332
rect 9355 22330 9411 22332
rect 9115 22278 9161 22330
rect 9161 22278 9171 22330
rect 9195 22278 9225 22330
rect 9225 22278 9237 22330
rect 9237 22278 9251 22330
rect 9275 22278 9289 22330
rect 9289 22278 9301 22330
rect 9301 22278 9331 22330
rect 9355 22278 9365 22330
rect 9365 22278 9411 22330
rect 9115 22276 9171 22278
rect 9195 22276 9251 22278
rect 9275 22276 9331 22278
rect 9355 22276 9411 22278
rect 10046 22500 10102 22536
rect 10046 22480 10048 22500
rect 10048 22480 10100 22500
rect 10100 22480 10102 22500
rect 9115 21242 9171 21244
rect 9195 21242 9251 21244
rect 9275 21242 9331 21244
rect 9355 21242 9411 21244
rect 9115 21190 9161 21242
rect 9161 21190 9171 21242
rect 9195 21190 9225 21242
rect 9225 21190 9237 21242
rect 9237 21190 9251 21242
rect 9275 21190 9289 21242
rect 9289 21190 9301 21242
rect 9301 21190 9331 21242
rect 9355 21190 9365 21242
rect 9365 21190 9411 21242
rect 9115 21188 9171 21190
rect 9195 21188 9251 21190
rect 9275 21188 9331 21190
rect 9355 21188 9411 21190
rect 9115 20154 9171 20156
rect 9195 20154 9251 20156
rect 9275 20154 9331 20156
rect 9355 20154 9411 20156
rect 9115 20102 9161 20154
rect 9161 20102 9171 20154
rect 9195 20102 9225 20154
rect 9225 20102 9237 20154
rect 9237 20102 9251 20154
rect 9275 20102 9289 20154
rect 9289 20102 9301 20154
rect 9301 20102 9331 20154
rect 9355 20102 9365 20154
rect 9365 20102 9411 20154
rect 9115 20100 9171 20102
rect 9195 20100 9251 20102
rect 9275 20100 9331 20102
rect 9355 20100 9411 20102
rect 9115 19066 9171 19068
rect 9195 19066 9251 19068
rect 9275 19066 9331 19068
rect 9355 19066 9411 19068
rect 9115 19014 9161 19066
rect 9161 19014 9171 19066
rect 9195 19014 9225 19066
rect 9225 19014 9237 19066
rect 9237 19014 9251 19066
rect 9275 19014 9289 19066
rect 9289 19014 9301 19066
rect 9301 19014 9331 19066
rect 9355 19014 9365 19066
rect 9365 19014 9411 19066
rect 9115 19012 9171 19014
rect 9195 19012 9251 19014
rect 9275 19012 9331 19014
rect 9355 19012 9411 19014
rect 10046 21836 10048 21856
rect 10048 21836 10100 21856
rect 10100 21836 10102 21856
rect 10046 21800 10102 21836
rect 10046 20984 10102 21040
rect 10046 20324 10102 20360
rect 10046 20304 10048 20324
rect 10048 20304 10100 20324
rect 10100 20304 10102 20324
rect 10046 19488 10102 19544
rect 9115 17978 9171 17980
rect 9195 17978 9251 17980
rect 9275 17978 9331 17980
rect 9355 17978 9411 17980
rect 9115 17926 9161 17978
rect 9161 17926 9171 17978
rect 9195 17926 9225 17978
rect 9225 17926 9237 17978
rect 9237 17926 9251 17978
rect 9275 17926 9289 17978
rect 9289 17926 9301 17978
rect 9301 17926 9331 17978
rect 9355 17926 9365 17978
rect 9365 17926 9411 17978
rect 9115 17924 9171 17926
rect 9195 17924 9251 17926
rect 9275 17924 9331 17926
rect 9355 17924 9411 17926
rect 9115 16890 9171 16892
rect 9195 16890 9251 16892
rect 9275 16890 9331 16892
rect 9355 16890 9411 16892
rect 9115 16838 9161 16890
rect 9161 16838 9171 16890
rect 9195 16838 9225 16890
rect 9225 16838 9237 16890
rect 9237 16838 9251 16890
rect 9275 16838 9289 16890
rect 9289 16838 9301 16890
rect 9301 16838 9331 16890
rect 9355 16838 9365 16890
rect 9365 16838 9411 16890
rect 9115 16836 9171 16838
rect 9195 16836 9251 16838
rect 9275 16836 9331 16838
rect 9355 16836 9411 16838
rect 9115 15802 9171 15804
rect 9195 15802 9251 15804
rect 9275 15802 9331 15804
rect 9355 15802 9411 15804
rect 9115 15750 9161 15802
rect 9161 15750 9171 15802
rect 9195 15750 9225 15802
rect 9225 15750 9237 15802
rect 9237 15750 9251 15802
rect 9275 15750 9289 15802
rect 9289 15750 9301 15802
rect 9301 15750 9331 15802
rect 9355 15750 9365 15802
rect 9365 15750 9411 15802
rect 9115 15748 9171 15750
rect 9195 15748 9251 15750
rect 9275 15748 9331 15750
rect 9355 15748 9411 15750
rect 9115 14714 9171 14716
rect 9195 14714 9251 14716
rect 9275 14714 9331 14716
rect 9355 14714 9411 14716
rect 9115 14662 9161 14714
rect 9161 14662 9171 14714
rect 9195 14662 9225 14714
rect 9225 14662 9237 14714
rect 9237 14662 9251 14714
rect 9275 14662 9289 14714
rect 9289 14662 9301 14714
rect 9301 14662 9331 14714
rect 9355 14662 9365 14714
rect 9365 14662 9411 14714
rect 9115 14660 9171 14662
rect 9195 14660 9251 14662
rect 9275 14660 9331 14662
rect 9355 14660 9411 14662
rect 10046 18672 10102 18728
rect 10046 18028 10048 18048
rect 10048 18028 10100 18048
rect 10100 18028 10102 18048
rect 10046 17992 10102 18028
rect 10046 17176 10102 17232
rect 10046 16396 10048 16416
rect 10048 16396 10100 16416
rect 10100 16396 10102 16416
rect 10046 16360 10102 16396
rect 10046 15680 10102 15736
rect 10046 14884 10102 14920
rect 10046 14864 10048 14884
rect 10048 14864 10100 14884
rect 10100 14864 10102 14884
rect 10046 14048 10102 14104
rect 9115 13626 9171 13628
rect 9195 13626 9251 13628
rect 9275 13626 9331 13628
rect 9355 13626 9411 13628
rect 9115 13574 9161 13626
rect 9161 13574 9171 13626
rect 9195 13574 9225 13626
rect 9225 13574 9237 13626
rect 9237 13574 9251 13626
rect 9275 13574 9289 13626
rect 9289 13574 9301 13626
rect 9301 13574 9331 13626
rect 9355 13574 9365 13626
rect 9365 13574 9411 13626
rect 9115 13572 9171 13574
rect 9195 13572 9251 13574
rect 9275 13572 9331 13574
rect 9355 13572 9411 13574
rect 10046 13368 10102 13424
rect 9115 12538 9171 12540
rect 9195 12538 9251 12540
rect 9275 12538 9331 12540
rect 9355 12538 9411 12540
rect 9115 12486 9161 12538
rect 9161 12486 9171 12538
rect 9195 12486 9225 12538
rect 9225 12486 9237 12538
rect 9237 12486 9251 12538
rect 9275 12486 9289 12538
rect 9289 12486 9301 12538
rect 9301 12486 9331 12538
rect 9355 12486 9365 12538
rect 9365 12486 9411 12538
rect 9115 12484 9171 12486
rect 9195 12484 9251 12486
rect 9275 12484 9331 12486
rect 9355 12484 9411 12486
rect 10046 12588 10048 12608
rect 10048 12588 10100 12608
rect 10100 12588 10102 12608
rect 10046 12552 10102 12588
rect 10046 11736 10102 11792
rect 9115 11450 9171 11452
rect 9195 11450 9251 11452
rect 9275 11450 9331 11452
rect 9355 11450 9411 11452
rect 9115 11398 9161 11450
rect 9161 11398 9171 11450
rect 9195 11398 9225 11450
rect 9225 11398 9237 11450
rect 9237 11398 9251 11450
rect 9275 11398 9289 11450
rect 9289 11398 9301 11450
rect 9301 11398 9331 11450
rect 9355 11398 9365 11450
rect 9365 11398 9411 11450
rect 9115 11396 9171 11398
rect 9195 11396 9251 11398
rect 9275 11396 9331 11398
rect 9355 11396 9411 11398
rect 10046 11056 10102 11112
rect 9115 10362 9171 10364
rect 9195 10362 9251 10364
rect 9275 10362 9331 10364
rect 9355 10362 9411 10364
rect 9115 10310 9161 10362
rect 9161 10310 9171 10362
rect 9195 10310 9225 10362
rect 9225 10310 9237 10362
rect 9237 10310 9251 10362
rect 9275 10310 9289 10362
rect 9289 10310 9301 10362
rect 9301 10310 9331 10362
rect 9355 10310 9365 10362
rect 9365 10310 9411 10362
rect 9115 10308 9171 10310
rect 9195 10308 9251 10310
rect 9275 10308 9331 10310
rect 9355 10308 9411 10310
rect 10046 10240 10102 10296
rect 9115 9274 9171 9276
rect 9195 9274 9251 9276
rect 9275 9274 9331 9276
rect 9355 9274 9411 9276
rect 9115 9222 9161 9274
rect 9161 9222 9171 9274
rect 9195 9222 9225 9274
rect 9225 9222 9237 9274
rect 9237 9222 9251 9274
rect 9275 9222 9289 9274
rect 9289 9222 9301 9274
rect 9301 9222 9331 9274
rect 9355 9222 9365 9274
rect 9365 9222 9411 9274
rect 9115 9220 9171 9222
rect 9195 9220 9251 9222
rect 9275 9220 9331 9222
rect 9355 9220 9411 9222
rect 10046 9444 10102 9480
rect 10046 9424 10048 9444
rect 10048 9424 10100 9444
rect 10100 9424 10102 9444
rect 10046 8780 10048 8800
rect 10048 8780 10100 8800
rect 10100 8780 10102 8800
rect 10046 8744 10102 8780
rect 9115 8186 9171 8188
rect 9195 8186 9251 8188
rect 9275 8186 9331 8188
rect 9355 8186 9411 8188
rect 9115 8134 9161 8186
rect 9161 8134 9171 8186
rect 9195 8134 9225 8186
rect 9225 8134 9237 8186
rect 9237 8134 9251 8186
rect 9275 8134 9289 8186
rect 9289 8134 9301 8186
rect 9301 8134 9331 8186
rect 9355 8134 9365 8186
rect 9365 8134 9411 8186
rect 9115 8132 9171 8134
rect 9195 8132 9251 8134
rect 9275 8132 9331 8134
rect 9355 8132 9411 8134
rect 10046 7928 10102 7984
rect 10046 7148 10048 7168
rect 10048 7148 10100 7168
rect 10100 7148 10102 7168
rect 9115 7098 9171 7100
rect 9195 7098 9251 7100
rect 9275 7098 9331 7100
rect 9355 7098 9411 7100
rect 9115 7046 9161 7098
rect 9161 7046 9171 7098
rect 9195 7046 9225 7098
rect 9225 7046 9237 7098
rect 9237 7046 9251 7098
rect 9275 7046 9289 7098
rect 9289 7046 9301 7098
rect 9301 7046 9331 7098
rect 9355 7046 9365 7098
rect 9365 7046 9411 7098
rect 9115 7044 9171 7046
rect 9195 7044 9251 7046
rect 9275 7044 9331 7046
rect 9355 7044 9411 7046
rect 7483 6554 7539 6556
rect 7563 6554 7619 6556
rect 7643 6554 7699 6556
rect 7723 6554 7779 6556
rect 7483 6502 7529 6554
rect 7529 6502 7539 6554
rect 7563 6502 7593 6554
rect 7593 6502 7605 6554
rect 7605 6502 7619 6554
rect 7643 6502 7657 6554
rect 7657 6502 7669 6554
rect 7669 6502 7699 6554
rect 7723 6502 7733 6554
rect 7733 6502 7779 6554
rect 7483 6500 7539 6502
rect 7563 6500 7619 6502
rect 7643 6500 7699 6502
rect 7723 6500 7779 6502
rect 5851 6010 5907 6012
rect 5931 6010 5987 6012
rect 6011 6010 6067 6012
rect 6091 6010 6147 6012
rect 5851 5958 5897 6010
rect 5897 5958 5907 6010
rect 5931 5958 5961 6010
rect 5961 5958 5973 6010
rect 5973 5958 5987 6010
rect 6011 5958 6025 6010
rect 6025 5958 6037 6010
rect 6037 5958 6067 6010
rect 6091 5958 6101 6010
rect 6101 5958 6147 6010
rect 5851 5956 5907 5958
rect 5931 5956 5987 5958
rect 6011 5956 6067 5958
rect 6091 5956 6147 5958
rect 7483 5466 7539 5468
rect 7563 5466 7619 5468
rect 7643 5466 7699 5468
rect 7723 5466 7779 5468
rect 7483 5414 7529 5466
rect 7529 5414 7539 5466
rect 7563 5414 7593 5466
rect 7593 5414 7605 5466
rect 7605 5414 7619 5466
rect 7643 5414 7657 5466
rect 7657 5414 7669 5466
rect 7669 5414 7699 5466
rect 7723 5414 7733 5466
rect 7733 5414 7779 5466
rect 7483 5412 7539 5414
rect 7563 5412 7619 5414
rect 7643 5412 7699 5414
rect 7723 5412 7779 5414
rect 5851 4922 5907 4924
rect 5931 4922 5987 4924
rect 6011 4922 6067 4924
rect 6091 4922 6147 4924
rect 5851 4870 5897 4922
rect 5897 4870 5907 4922
rect 5931 4870 5961 4922
rect 5961 4870 5973 4922
rect 5973 4870 5987 4922
rect 6011 4870 6025 4922
rect 6025 4870 6037 4922
rect 6037 4870 6067 4922
rect 6091 4870 6101 4922
rect 6101 4870 6147 4922
rect 5851 4868 5907 4870
rect 5931 4868 5987 4870
rect 6011 4868 6067 4870
rect 6091 4868 6147 4870
rect 7483 4378 7539 4380
rect 7563 4378 7619 4380
rect 7643 4378 7699 4380
rect 7723 4378 7779 4380
rect 7483 4326 7529 4378
rect 7529 4326 7539 4378
rect 7563 4326 7593 4378
rect 7593 4326 7605 4378
rect 7605 4326 7619 4378
rect 7643 4326 7657 4378
rect 7657 4326 7669 4378
rect 7669 4326 7699 4378
rect 7723 4326 7733 4378
rect 7733 4326 7779 4378
rect 7483 4324 7539 4326
rect 7563 4324 7619 4326
rect 7643 4324 7699 4326
rect 7723 4324 7779 4326
rect 5851 3834 5907 3836
rect 5931 3834 5987 3836
rect 6011 3834 6067 3836
rect 6091 3834 6147 3836
rect 5851 3782 5897 3834
rect 5897 3782 5907 3834
rect 5931 3782 5961 3834
rect 5961 3782 5973 3834
rect 5973 3782 5987 3834
rect 6011 3782 6025 3834
rect 6025 3782 6037 3834
rect 6037 3782 6067 3834
rect 6091 3782 6101 3834
rect 6101 3782 6147 3834
rect 5851 3780 5907 3782
rect 5931 3780 5987 3782
rect 6011 3780 6067 3782
rect 6091 3780 6147 3782
rect 9115 6010 9171 6012
rect 9195 6010 9251 6012
rect 9275 6010 9331 6012
rect 9355 6010 9411 6012
rect 9115 5958 9161 6010
rect 9161 5958 9171 6010
rect 9195 5958 9225 6010
rect 9225 5958 9237 6010
rect 9237 5958 9251 6010
rect 9275 5958 9289 6010
rect 9289 5958 9301 6010
rect 9301 5958 9331 6010
rect 9355 5958 9365 6010
rect 9365 5958 9411 6010
rect 9115 5956 9171 5958
rect 9195 5956 9251 5958
rect 9275 5956 9331 5958
rect 9355 5956 9411 5958
rect 10046 7112 10102 7148
rect 10046 6432 10102 6488
rect 10046 5616 10102 5672
rect 9115 4922 9171 4924
rect 9195 4922 9251 4924
rect 9275 4922 9331 4924
rect 9355 4922 9411 4924
rect 9115 4870 9161 4922
rect 9161 4870 9171 4922
rect 9195 4870 9225 4922
rect 9225 4870 9237 4922
rect 9237 4870 9251 4922
rect 9275 4870 9289 4922
rect 9289 4870 9301 4922
rect 9301 4870 9331 4922
rect 9355 4870 9365 4922
rect 9365 4870 9411 4922
rect 9115 4868 9171 4870
rect 9195 4868 9251 4870
rect 9275 4868 9331 4870
rect 9355 4868 9411 4870
rect 10046 4800 10102 4856
rect 7483 3290 7539 3292
rect 7563 3290 7619 3292
rect 7643 3290 7699 3292
rect 7723 3290 7779 3292
rect 7483 3238 7529 3290
rect 7529 3238 7539 3290
rect 7563 3238 7593 3290
rect 7593 3238 7605 3290
rect 7605 3238 7619 3290
rect 7643 3238 7657 3290
rect 7657 3238 7669 3290
rect 7669 3238 7699 3290
rect 7723 3238 7733 3290
rect 7733 3238 7779 3290
rect 7483 3236 7539 3238
rect 7563 3236 7619 3238
rect 7643 3236 7699 3238
rect 7723 3236 7779 3238
rect 9115 3834 9171 3836
rect 9195 3834 9251 3836
rect 9275 3834 9331 3836
rect 9355 3834 9411 3836
rect 9115 3782 9161 3834
rect 9161 3782 9171 3834
rect 9195 3782 9225 3834
rect 9225 3782 9237 3834
rect 9237 3782 9251 3834
rect 9275 3782 9289 3834
rect 9289 3782 9301 3834
rect 9301 3782 9331 3834
rect 9355 3782 9365 3834
rect 9365 3782 9411 3834
rect 9115 3780 9171 3782
rect 9195 3780 9251 3782
rect 9275 3780 9331 3782
rect 9355 3780 9411 3782
rect 10046 4120 10102 4176
rect 10046 3340 10048 3360
rect 10048 3340 10100 3360
rect 10100 3340 10102 3360
rect 10046 3304 10102 3340
rect 5851 2746 5907 2748
rect 5931 2746 5987 2748
rect 6011 2746 6067 2748
rect 6091 2746 6147 2748
rect 5851 2694 5897 2746
rect 5897 2694 5907 2746
rect 5931 2694 5961 2746
rect 5961 2694 5973 2746
rect 5973 2694 5987 2746
rect 6011 2694 6025 2746
rect 6025 2694 6037 2746
rect 6037 2694 6067 2746
rect 6091 2694 6101 2746
rect 6101 2694 6147 2746
rect 5851 2692 5907 2694
rect 5931 2692 5987 2694
rect 6011 2692 6067 2694
rect 6091 2692 6147 2694
rect 9115 2746 9171 2748
rect 9195 2746 9251 2748
rect 9275 2746 9331 2748
rect 9355 2746 9411 2748
rect 9115 2694 9161 2746
rect 9161 2694 9171 2746
rect 9195 2694 9225 2746
rect 9225 2694 9237 2746
rect 9237 2694 9251 2746
rect 9275 2694 9289 2746
rect 9289 2694 9301 2746
rect 9301 2694 9331 2746
rect 9355 2694 9365 2746
rect 9365 2694 9411 2746
rect 9115 2692 9171 2694
rect 9195 2692 9251 2694
rect 9275 2692 9331 2694
rect 9355 2692 9411 2694
rect 3606 2216 3662 2272
rect 4219 2202 4275 2204
rect 4299 2202 4355 2204
rect 4379 2202 4435 2204
rect 4459 2202 4515 2204
rect 4219 2150 4265 2202
rect 4265 2150 4275 2202
rect 4299 2150 4329 2202
rect 4329 2150 4341 2202
rect 4341 2150 4355 2202
rect 4379 2150 4393 2202
rect 4393 2150 4405 2202
rect 4405 2150 4435 2202
rect 4459 2150 4469 2202
rect 4469 2150 4515 2202
rect 4219 2148 4275 2150
rect 4299 2148 4355 2150
rect 4379 2148 4435 2150
rect 4459 2148 4515 2150
rect 3974 1808 4030 1864
rect 2870 1400 2926 1456
rect 2870 1028 2872 1048
rect 2872 1028 2924 1048
rect 2924 1028 2926 1048
rect 2870 992 2926 1028
rect 2778 584 2834 640
rect 2778 176 2834 232
rect 7483 2202 7539 2204
rect 7563 2202 7619 2204
rect 7643 2202 7699 2204
rect 7723 2202 7779 2204
rect 7483 2150 7529 2202
rect 7529 2150 7539 2202
rect 7563 2150 7593 2202
rect 7593 2150 7605 2202
rect 7605 2150 7619 2202
rect 7643 2150 7657 2202
rect 7657 2150 7669 2202
rect 7669 2150 7699 2202
rect 7723 2150 7733 2202
rect 7733 2150 7779 2202
rect 7483 2148 7539 2150
rect 7563 2148 7619 2150
rect 7643 2148 7699 2150
rect 7723 2148 7779 2150
rect 10046 2488 10102 2544
rect 9494 1808 9550 1864
rect 10046 992 10102 1048
rect 9310 312 9366 368
<< metal3 >>
rect 0 79658 800 79688
rect 2957 79658 3023 79661
rect 0 79656 3023 79658
rect 0 79600 2962 79656
rect 3018 79600 3023 79656
rect 0 79598 3023 79600
rect 0 79568 800 79598
rect 2957 79595 3023 79598
rect 10041 79522 10107 79525
rect 11200 79522 12000 79552
rect 10041 79520 12000 79522
rect 10041 79464 10046 79520
rect 10102 79464 12000 79520
rect 10041 79462 12000 79464
rect 10041 79459 10107 79462
rect 11200 79432 12000 79462
rect 0 79250 800 79280
rect 1393 79250 1459 79253
rect 0 79248 1459 79250
rect 0 79192 1398 79248
rect 1454 79192 1459 79248
rect 0 79190 1459 79192
rect 0 79160 800 79190
rect 1393 79187 1459 79190
rect 0 78842 800 78872
rect 2773 78842 2839 78845
rect 0 78840 2839 78842
rect 0 78784 2778 78840
rect 2834 78784 2839 78840
rect 0 78782 2839 78784
rect 0 78752 800 78782
rect 2773 78779 2839 78782
rect 10961 78706 11027 78709
rect 11200 78706 12000 78736
rect 10961 78704 12000 78706
rect 10961 78648 10966 78704
rect 11022 78648 12000 78704
rect 10961 78646 12000 78648
rect 10961 78643 11027 78646
rect 11200 78616 12000 78646
rect 0 78434 800 78464
rect 3509 78434 3575 78437
rect 0 78432 3575 78434
rect 0 78376 3514 78432
rect 3570 78376 3575 78432
rect 0 78374 3575 78376
rect 0 78344 800 78374
rect 3509 78371 3575 78374
rect 0 78026 800 78056
rect 4061 78026 4127 78029
rect 0 78024 4127 78026
rect 0 77968 4066 78024
rect 4122 77968 4127 78024
rect 0 77966 4127 77968
rect 0 77936 800 77966
rect 4061 77963 4127 77966
rect 9489 78026 9555 78029
rect 11200 78026 12000 78056
rect 9489 78024 12000 78026
rect 9489 77968 9494 78024
rect 9550 77968 12000 78024
rect 9489 77966 12000 77968
rect 9489 77963 9555 77966
rect 11200 77936 12000 77966
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5839 77824 6159 77825
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 77759 6159 77760
rect 9103 77824 9423 77825
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 77759 9423 77760
rect 0 77618 800 77648
rect 3417 77618 3483 77621
rect 0 77616 3483 77618
rect 0 77560 3422 77616
rect 3478 77560 3483 77616
rect 0 77558 3483 77560
rect 0 77528 800 77558
rect 3417 77555 3483 77558
rect 4207 77280 4527 77281
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 77215 4527 77216
rect 7471 77280 7791 77281
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 77215 7791 77216
rect 9397 77210 9463 77213
rect 11200 77210 12000 77240
rect 9397 77208 12000 77210
rect 9397 77152 9402 77208
rect 9458 77152 12000 77208
rect 9397 77150 12000 77152
rect 9397 77147 9463 77150
rect 11200 77120 12000 77150
rect 0 77074 800 77104
rect 3969 77074 4035 77077
rect 0 77072 4035 77074
rect 0 77016 3974 77072
rect 4030 77016 4035 77072
rect 0 77014 4035 77016
rect 0 76984 800 77014
rect 3969 77011 4035 77014
rect 2576 76736 2896 76737
rect 0 76666 800 76696
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5839 76736 6159 76737
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 76671 6159 76672
rect 9103 76736 9423 76737
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 76671 9423 76672
rect 0 76606 1778 76666
rect 0 76576 800 76606
rect 1718 76530 1778 76606
rect 3325 76530 3391 76533
rect 1718 76528 3391 76530
rect 1718 76472 3330 76528
rect 3386 76472 3391 76528
rect 1718 76470 3391 76472
rect 3325 76467 3391 76470
rect 10133 76394 10199 76397
rect 11200 76394 12000 76424
rect 10133 76392 12000 76394
rect 10133 76336 10138 76392
rect 10194 76336 12000 76392
rect 10133 76334 12000 76336
rect 10133 76331 10199 76334
rect 11200 76304 12000 76334
rect 0 76258 800 76288
rect 2957 76258 3023 76261
rect 0 76256 3023 76258
rect 0 76200 2962 76256
rect 3018 76200 3023 76256
rect 0 76198 3023 76200
rect 0 76168 800 76198
rect 2957 76195 3023 76198
rect 4207 76192 4527 76193
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 76127 4527 76128
rect 7471 76192 7791 76193
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 76127 7791 76128
rect 0 75850 800 75880
rect 3141 75850 3207 75853
rect 0 75848 3207 75850
rect 0 75792 3146 75848
rect 3202 75792 3207 75848
rect 0 75790 3207 75792
rect 0 75760 800 75790
rect 3141 75787 3207 75790
rect 10225 75714 10291 75717
rect 11200 75714 12000 75744
rect 10225 75712 12000 75714
rect 10225 75656 10230 75712
rect 10286 75656 12000 75712
rect 10225 75654 12000 75656
rect 10225 75651 10291 75654
rect 2576 75648 2896 75649
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5839 75648 6159 75649
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 75583 6159 75584
rect 9103 75648 9423 75649
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 11200 75624 12000 75654
rect 9103 75583 9423 75584
rect 0 75442 800 75472
rect 3601 75442 3667 75445
rect 0 75440 3667 75442
rect 0 75384 3606 75440
rect 3662 75384 3667 75440
rect 0 75382 3667 75384
rect 0 75352 800 75382
rect 3601 75379 3667 75382
rect 4207 75104 4527 75105
rect 0 75034 800 75064
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 75039 4527 75040
rect 7471 75104 7791 75105
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 75039 7791 75040
rect 3141 75034 3207 75037
rect 0 75032 3207 75034
rect 0 74976 3146 75032
rect 3202 74976 3207 75032
rect 0 74974 3207 74976
rect 0 74944 800 74974
rect 3141 74971 3207 74974
rect 10133 74898 10199 74901
rect 11200 74898 12000 74928
rect 10133 74896 12000 74898
rect 10133 74840 10138 74896
rect 10194 74840 12000 74896
rect 10133 74838 12000 74840
rect 10133 74835 10199 74838
rect 11200 74808 12000 74838
rect 2576 74560 2896 74561
rect 0 74490 800 74520
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5839 74560 6159 74561
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 74495 6159 74496
rect 9103 74560 9423 74561
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 74495 9423 74496
rect 1485 74490 1551 74493
rect 0 74488 1551 74490
rect 0 74432 1490 74488
rect 1546 74432 1551 74488
rect 0 74430 1551 74432
rect 0 74400 800 74430
rect 1485 74427 1551 74430
rect 1393 74354 1459 74357
rect 982 74352 1459 74354
rect 982 74296 1398 74352
rect 1454 74296 1459 74352
rect 982 74294 1459 74296
rect 0 74082 800 74112
rect 982 74082 1042 74294
rect 1393 74291 1459 74294
rect 0 74022 1042 74082
rect 10133 74082 10199 74085
rect 11200 74082 12000 74112
rect 10133 74080 12000 74082
rect 10133 74024 10138 74080
rect 10194 74024 12000 74080
rect 10133 74022 12000 74024
rect 0 73992 800 74022
rect 10133 74019 10199 74022
rect 4207 74016 4527 74017
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 73951 4527 73952
rect 7471 74016 7791 74017
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 11200 73992 12000 74022
rect 7471 73951 7791 73952
rect 0 73674 800 73704
rect 2773 73674 2839 73677
rect 0 73672 2839 73674
rect 0 73616 2778 73672
rect 2834 73616 2839 73672
rect 0 73614 2839 73616
rect 0 73584 800 73614
rect 2773 73611 2839 73614
rect 2576 73472 2896 73473
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5839 73472 6159 73473
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 73407 6159 73408
rect 9103 73472 9423 73473
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 73407 9423 73408
rect 10133 73402 10199 73405
rect 11200 73402 12000 73432
rect 10133 73400 12000 73402
rect 10133 73344 10138 73400
rect 10194 73344 12000 73400
rect 10133 73342 12000 73344
rect 10133 73339 10199 73342
rect 11200 73312 12000 73342
rect 0 73266 800 73296
rect 1393 73266 1459 73269
rect 0 73264 1459 73266
rect 0 73208 1398 73264
rect 1454 73208 1459 73264
rect 0 73206 1459 73208
rect 0 73176 800 73206
rect 1393 73203 1459 73206
rect 4207 72928 4527 72929
rect 0 72858 800 72888
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 72863 4527 72864
rect 7471 72928 7791 72929
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 72863 7791 72864
rect 2773 72858 2839 72861
rect 0 72856 2839 72858
rect 0 72800 2778 72856
rect 2834 72800 2839 72856
rect 0 72798 2839 72800
rect 0 72768 800 72798
rect 2773 72795 2839 72798
rect 10133 72586 10199 72589
rect 11200 72586 12000 72616
rect 10133 72584 12000 72586
rect 10133 72528 10138 72584
rect 10194 72528 12000 72584
rect 10133 72526 12000 72528
rect 10133 72523 10199 72526
rect 11200 72496 12000 72526
rect 0 72450 800 72480
rect 2037 72450 2103 72453
rect 0 72448 2103 72450
rect 0 72392 2042 72448
rect 2098 72392 2103 72448
rect 0 72390 2103 72392
rect 0 72360 800 72390
rect 2037 72387 2103 72390
rect 2576 72384 2896 72385
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5839 72384 6159 72385
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 72319 6159 72320
rect 9103 72384 9423 72385
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 72319 9423 72320
rect 0 71906 800 71936
rect 1393 71906 1459 71909
rect 0 71904 1459 71906
rect 0 71848 1398 71904
rect 1454 71848 1459 71904
rect 0 71846 1459 71848
rect 0 71816 800 71846
rect 1393 71843 1459 71846
rect 4207 71840 4527 71841
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 71775 4527 71776
rect 7471 71840 7791 71841
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 71775 7791 71776
rect 10133 71770 10199 71773
rect 11200 71770 12000 71800
rect 10133 71768 12000 71770
rect 10133 71712 10138 71768
rect 10194 71712 12000 71768
rect 10133 71710 12000 71712
rect 10133 71707 10199 71710
rect 11200 71680 12000 71710
rect 0 71498 800 71528
rect 2221 71498 2287 71501
rect 0 71496 2287 71498
rect 0 71440 2226 71496
rect 2282 71440 2287 71496
rect 0 71438 2287 71440
rect 0 71408 800 71438
rect 2221 71435 2287 71438
rect 2576 71296 2896 71297
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5839 71296 6159 71297
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 71231 6159 71232
rect 9103 71296 9423 71297
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 71231 9423 71232
rect 0 71090 800 71120
rect 1209 71090 1275 71093
rect 0 71088 1275 71090
rect 0 71032 1214 71088
rect 1270 71032 1275 71088
rect 0 71030 1275 71032
rect 0 71000 800 71030
rect 1209 71027 1275 71030
rect 10133 71090 10199 71093
rect 11200 71090 12000 71120
rect 10133 71088 12000 71090
rect 10133 71032 10138 71088
rect 10194 71032 12000 71088
rect 10133 71030 12000 71032
rect 10133 71027 10199 71030
rect 11200 71000 12000 71030
rect 4207 70752 4527 70753
rect 0 70682 800 70712
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 70687 4527 70688
rect 7471 70752 7791 70753
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 70687 7791 70688
rect 1301 70682 1367 70685
rect 0 70680 1367 70682
rect 0 70624 1306 70680
rect 1362 70624 1367 70680
rect 0 70622 1367 70624
rect 0 70592 800 70622
rect 1301 70619 1367 70622
rect 0 70274 800 70304
rect 1393 70274 1459 70277
rect 0 70272 1459 70274
rect 0 70216 1398 70272
rect 1454 70216 1459 70272
rect 0 70214 1459 70216
rect 0 70184 800 70214
rect 1393 70211 1459 70214
rect 10133 70274 10199 70277
rect 11200 70274 12000 70304
rect 10133 70272 12000 70274
rect 10133 70216 10138 70272
rect 10194 70216 12000 70272
rect 10133 70214 12000 70216
rect 10133 70211 10199 70214
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5839 70208 6159 70209
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 70143 6159 70144
rect 9103 70208 9423 70209
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 11200 70184 12000 70214
rect 9103 70143 9423 70144
rect 0 69866 800 69896
rect 2957 69866 3023 69869
rect 0 69864 3023 69866
rect 0 69808 2962 69864
rect 3018 69808 3023 69864
rect 0 69806 3023 69808
rect 0 69776 800 69806
rect 2957 69803 3023 69806
rect 4207 69664 4527 69665
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 69599 4527 69600
rect 7471 69664 7791 69665
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 69599 7791 69600
rect 10133 69458 10199 69461
rect 11200 69458 12000 69488
rect 10133 69456 12000 69458
rect 10133 69400 10138 69456
rect 10194 69400 12000 69456
rect 10133 69398 12000 69400
rect 10133 69395 10199 69398
rect 11200 69368 12000 69398
rect 0 69322 800 69352
rect 3325 69322 3391 69325
rect 0 69320 3391 69322
rect 0 69264 3330 69320
rect 3386 69264 3391 69320
rect 0 69262 3391 69264
rect 0 69232 800 69262
rect 3325 69259 3391 69262
rect 2576 69120 2896 69121
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5839 69120 6159 69121
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 69055 6159 69056
rect 9103 69120 9423 69121
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 69055 9423 69056
rect 0 68914 800 68944
rect 3049 68914 3115 68917
rect 0 68912 3115 68914
rect 0 68856 3054 68912
rect 3110 68856 3115 68912
rect 0 68854 3115 68856
rect 0 68824 800 68854
rect 3049 68851 3115 68854
rect 1301 68778 1367 68781
rect 2865 68778 2931 68781
rect 1301 68776 2931 68778
rect 1301 68720 1306 68776
rect 1362 68720 2870 68776
rect 2926 68720 2931 68776
rect 1301 68718 2931 68720
rect 1301 68715 1367 68718
rect 2865 68715 2931 68718
rect 10133 68778 10199 68781
rect 11200 68778 12000 68808
rect 10133 68776 12000 68778
rect 10133 68720 10138 68776
rect 10194 68720 12000 68776
rect 10133 68718 12000 68720
rect 10133 68715 10199 68718
rect 11200 68688 12000 68718
rect 4207 68576 4527 68577
rect 0 68506 800 68536
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 68511 4527 68512
rect 7471 68576 7791 68577
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 68511 7791 68512
rect 2957 68506 3023 68509
rect 0 68504 3023 68506
rect 0 68448 2962 68504
rect 3018 68448 3023 68504
rect 0 68446 3023 68448
rect 0 68416 800 68446
rect 2957 68443 3023 68446
rect 0 68098 800 68128
rect 1393 68098 1459 68101
rect 0 68096 1459 68098
rect 0 68040 1398 68096
rect 1454 68040 1459 68096
rect 0 68038 1459 68040
rect 0 68008 800 68038
rect 1393 68035 1459 68038
rect 2576 68032 2896 68033
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5839 68032 6159 68033
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 67967 6159 67968
rect 9103 68032 9423 68033
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 67967 9423 67968
rect 10133 67962 10199 67965
rect 11200 67962 12000 67992
rect 10133 67960 12000 67962
rect 10133 67904 10138 67960
rect 10194 67904 12000 67960
rect 10133 67902 12000 67904
rect 10133 67899 10199 67902
rect 11200 67872 12000 67902
rect 0 67690 800 67720
rect 1301 67690 1367 67693
rect 0 67688 1367 67690
rect 0 67632 1306 67688
rect 1362 67632 1367 67688
rect 0 67630 1367 67632
rect 0 67600 800 67630
rect 1301 67627 1367 67630
rect 4207 67488 4527 67489
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 67423 4527 67424
rect 7471 67488 7791 67489
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 67423 7791 67424
rect 0 67282 800 67312
rect 1393 67282 1459 67285
rect 0 67280 1459 67282
rect 0 67224 1398 67280
rect 1454 67224 1459 67280
rect 0 67222 1459 67224
rect 0 67192 800 67222
rect 1393 67219 1459 67222
rect 10133 67146 10199 67149
rect 11200 67146 12000 67176
rect 10133 67144 12000 67146
rect 10133 67088 10138 67144
rect 10194 67088 12000 67144
rect 10133 67086 12000 67088
rect 10133 67083 10199 67086
rect 11200 67056 12000 67086
rect 2576 66944 2896 66945
rect 0 66874 800 66904
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5839 66944 6159 66945
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 66879 6159 66880
rect 9103 66944 9423 66945
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 66879 9423 66880
rect 1393 66874 1459 66877
rect 0 66872 1459 66874
rect 0 66816 1398 66872
rect 1454 66816 1459 66872
rect 0 66814 1459 66816
rect 0 66784 800 66814
rect 1393 66811 1459 66814
rect 1761 66466 1827 66469
rect 2078 66466 2084 66468
rect 1761 66464 2084 66466
rect 1761 66408 1766 66464
rect 1822 66408 2084 66464
rect 1761 66406 2084 66408
rect 1761 66403 1827 66406
rect 2078 66404 2084 66406
rect 2148 66404 2154 66468
rect 10133 66466 10199 66469
rect 11200 66466 12000 66496
rect 10133 66464 12000 66466
rect 10133 66408 10138 66464
rect 10194 66408 12000 66464
rect 10133 66406 12000 66408
rect 10133 66403 10199 66406
rect 4207 66400 4527 66401
rect 0 66330 800 66360
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 66335 4527 66336
rect 7471 66400 7791 66401
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 11200 66376 12000 66406
rect 7471 66335 7791 66336
rect 1393 66330 1459 66333
rect 0 66328 1459 66330
rect 0 66272 1398 66328
rect 1454 66272 1459 66328
rect 0 66270 1459 66272
rect 0 66240 800 66270
rect 1393 66267 1459 66270
rect 1669 66194 1735 66197
rect 7189 66194 7255 66197
rect 1669 66192 7255 66194
rect 1669 66136 1674 66192
rect 1730 66136 7194 66192
rect 7250 66136 7255 66192
rect 1669 66134 7255 66136
rect 1669 66131 1735 66134
rect 7189 66131 7255 66134
rect 0 65922 800 65952
rect 1393 65922 1459 65925
rect 0 65920 1459 65922
rect 0 65864 1398 65920
rect 1454 65864 1459 65920
rect 0 65862 1459 65864
rect 0 65832 800 65862
rect 1393 65859 1459 65862
rect 2576 65856 2896 65857
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5839 65856 6159 65857
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 65791 6159 65792
rect 9103 65856 9423 65857
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 65791 9423 65792
rect 1761 65650 1827 65653
rect 5901 65650 5967 65653
rect 1761 65648 5967 65650
rect 1761 65592 1766 65648
rect 1822 65592 5906 65648
rect 5962 65592 5967 65648
rect 1761 65590 5967 65592
rect 1761 65587 1827 65590
rect 5901 65587 5967 65590
rect 10133 65650 10199 65653
rect 11200 65650 12000 65680
rect 10133 65648 12000 65650
rect 10133 65592 10138 65648
rect 10194 65592 12000 65648
rect 10133 65590 12000 65592
rect 10133 65587 10199 65590
rect 11200 65560 12000 65590
rect 0 65514 800 65544
rect 2957 65514 3023 65517
rect 0 65512 3023 65514
rect 0 65456 2962 65512
rect 3018 65456 3023 65512
rect 0 65454 3023 65456
rect 0 65424 800 65454
rect 2957 65451 3023 65454
rect 4207 65312 4527 65313
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 65247 4527 65248
rect 7471 65312 7791 65313
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 65247 7791 65248
rect 0 65106 800 65136
rect 3325 65106 3391 65109
rect 0 65104 3391 65106
rect 0 65048 3330 65104
rect 3386 65048 3391 65104
rect 0 65046 3391 65048
rect 0 65016 800 65046
rect 3325 65043 3391 65046
rect 1894 64908 1900 64972
rect 1964 64970 1970 64972
rect 2129 64970 2195 64973
rect 1964 64968 2195 64970
rect 1964 64912 2134 64968
rect 2190 64912 2195 64968
rect 1964 64910 2195 64912
rect 1964 64908 1970 64910
rect 2129 64907 2195 64910
rect 10133 64834 10199 64837
rect 11200 64834 12000 64864
rect 10133 64832 12000 64834
rect 10133 64776 10138 64832
rect 10194 64776 12000 64832
rect 10133 64774 12000 64776
rect 10133 64771 10199 64774
rect 2576 64768 2896 64769
rect 0 64698 800 64728
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 5839 64768 6159 64769
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 64703 6159 64704
rect 9103 64768 9423 64769
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 11200 64744 12000 64774
rect 9103 64703 9423 64704
rect 0 64638 1456 64698
rect 0 64608 800 64638
rect 1396 64562 1456 64638
rect 3877 64562 3943 64565
rect 1396 64560 3943 64562
rect 1396 64504 3882 64560
rect 3938 64504 3943 64560
rect 1396 64502 3943 64504
rect 3877 64499 3943 64502
rect 0 64290 800 64320
rect 2773 64290 2839 64293
rect 0 64288 2839 64290
rect 0 64232 2778 64288
rect 2834 64232 2839 64288
rect 0 64230 2839 64232
rect 0 64200 800 64230
rect 2773 64227 2839 64230
rect 4207 64224 4527 64225
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 64159 4527 64160
rect 7471 64224 7791 64225
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 64159 7791 64160
rect 10133 64154 10199 64157
rect 11200 64154 12000 64184
rect 10133 64152 12000 64154
rect 10133 64096 10138 64152
rect 10194 64096 12000 64152
rect 10133 64094 12000 64096
rect 10133 64091 10199 64094
rect 11200 64064 12000 64094
rect 0 63746 800 63776
rect 2221 63746 2287 63749
rect 0 63744 2287 63746
rect 0 63688 2226 63744
rect 2282 63688 2287 63744
rect 0 63686 2287 63688
rect 0 63656 800 63686
rect 2221 63683 2287 63686
rect 2576 63680 2896 63681
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5839 63680 6159 63681
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 63615 6159 63616
rect 9103 63680 9423 63681
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 63615 9423 63616
rect 0 63338 800 63368
rect 3049 63338 3115 63341
rect 0 63336 3115 63338
rect 0 63280 3054 63336
rect 3110 63280 3115 63336
rect 0 63278 3115 63280
rect 0 63248 800 63278
rect 3049 63275 3115 63278
rect 10133 63338 10199 63341
rect 11200 63338 12000 63368
rect 10133 63336 12000 63338
rect 10133 63280 10138 63336
rect 10194 63280 12000 63336
rect 10133 63278 12000 63280
rect 10133 63275 10199 63278
rect 11200 63248 12000 63278
rect 4207 63136 4527 63137
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 63071 4527 63072
rect 7471 63136 7791 63137
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 63071 7791 63072
rect 0 62930 800 62960
rect 2865 62930 2931 62933
rect 0 62928 2931 62930
rect 0 62872 2870 62928
rect 2926 62872 2931 62928
rect 0 62870 2931 62872
rect 0 62840 800 62870
rect 2865 62867 2931 62870
rect 2576 62592 2896 62593
rect 0 62522 800 62552
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5839 62592 6159 62593
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 62527 6159 62528
rect 9103 62592 9423 62593
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 62527 9423 62528
rect 1393 62522 1459 62525
rect 0 62520 1459 62522
rect 0 62464 1398 62520
rect 1454 62464 1459 62520
rect 0 62462 1459 62464
rect 0 62432 800 62462
rect 1393 62459 1459 62462
rect 10133 62522 10199 62525
rect 11200 62522 12000 62552
rect 10133 62520 12000 62522
rect 10133 62464 10138 62520
rect 10194 62464 12000 62520
rect 10133 62462 12000 62464
rect 10133 62459 10199 62462
rect 11200 62432 12000 62462
rect 0 62114 800 62144
rect 1485 62114 1551 62117
rect 0 62112 1551 62114
rect 0 62056 1490 62112
rect 1546 62056 1551 62112
rect 0 62054 1551 62056
rect 0 62024 800 62054
rect 1485 62051 1551 62054
rect 4207 62048 4527 62049
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 61983 4527 61984
rect 7471 62048 7791 62049
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 61983 7791 61984
rect 10133 61842 10199 61845
rect 11200 61842 12000 61872
rect 10133 61840 12000 61842
rect 10133 61784 10138 61840
rect 10194 61784 12000 61840
rect 10133 61782 12000 61784
rect 10133 61779 10199 61782
rect 11200 61752 12000 61782
rect 0 61706 800 61736
rect 1485 61706 1551 61709
rect 0 61704 1551 61706
rect 0 61648 1490 61704
rect 1546 61648 1551 61704
rect 0 61646 1551 61648
rect 0 61616 800 61646
rect 1485 61643 1551 61646
rect 2576 61504 2896 61505
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5839 61504 6159 61505
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 61439 6159 61440
rect 9103 61504 9423 61505
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 61439 9423 61440
rect 0 61162 800 61192
rect 1393 61162 1459 61165
rect 0 61160 1459 61162
rect 0 61104 1398 61160
rect 1454 61104 1459 61160
rect 0 61102 1459 61104
rect 0 61072 800 61102
rect 1393 61099 1459 61102
rect 10133 61026 10199 61029
rect 11200 61026 12000 61056
rect 10133 61024 12000 61026
rect 10133 60968 10138 61024
rect 10194 60968 12000 61024
rect 10133 60966 12000 60968
rect 10133 60963 10199 60966
rect 4207 60960 4527 60961
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 60895 4527 60896
rect 7471 60960 7791 60961
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 11200 60936 12000 60966
rect 7471 60895 7791 60896
rect 2262 60828 2268 60892
rect 2332 60890 2338 60892
rect 2497 60890 2563 60893
rect 2332 60888 2563 60890
rect 2332 60832 2502 60888
rect 2558 60832 2563 60888
rect 2332 60830 2563 60832
rect 2332 60828 2338 60830
rect 2497 60827 2563 60830
rect 0 60754 800 60784
rect 1485 60754 1551 60757
rect 0 60752 1551 60754
rect 0 60696 1490 60752
rect 1546 60696 1551 60752
rect 0 60694 1551 60696
rect 0 60664 800 60694
rect 1485 60691 1551 60694
rect 2078 60692 2084 60756
rect 2148 60754 2154 60756
rect 2497 60754 2563 60757
rect 2148 60752 2563 60754
rect 2148 60696 2502 60752
rect 2558 60696 2563 60752
rect 2148 60694 2563 60696
rect 2148 60692 2154 60694
rect 2497 60691 2563 60694
rect 2773 60618 2839 60621
rect 1396 60616 2839 60618
rect 1396 60560 2778 60616
rect 2834 60560 2839 60616
rect 1396 60558 2839 60560
rect 0 60346 800 60376
rect 1396 60346 1456 60558
rect 2773 60555 2839 60558
rect 2576 60416 2896 60417
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5839 60416 6159 60417
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 60351 6159 60352
rect 9103 60416 9423 60417
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 60351 9423 60352
rect 0 60286 1456 60346
rect 10133 60346 10199 60349
rect 11200 60346 12000 60376
rect 10133 60344 12000 60346
rect 10133 60288 10138 60344
rect 10194 60288 12000 60344
rect 10133 60286 12000 60288
rect 0 60256 800 60286
rect 10133 60283 10199 60286
rect 11200 60256 12000 60286
rect 2262 60148 2268 60212
rect 2332 60210 2338 60212
rect 2497 60210 2563 60213
rect 2332 60208 2563 60210
rect 2332 60152 2502 60208
rect 2558 60152 2563 60208
rect 2332 60150 2563 60152
rect 2332 60148 2338 60150
rect 2497 60147 2563 60150
rect 0 59938 800 59968
rect 1393 59938 1459 59941
rect 0 59936 1459 59938
rect 0 59880 1398 59936
rect 1454 59880 1459 59936
rect 0 59878 1459 59880
rect 0 59848 800 59878
rect 1393 59875 1459 59878
rect 4207 59872 4527 59873
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 59807 4527 59808
rect 7471 59872 7791 59873
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 59807 7791 59808
rect 1710 59604 1716 59668
rect 1780 59666 1786 59668
rect 2681 59666 2747 59669
rect 1780 59664 2747 59666
rect 1780 59608 2686 59664
rect 2742 59608 2747 59664
rect 1780 59606 2747 59608
rect 1780 59604 1786 59606
rect 2681 59603 2747 59606
rect 0 59530 800 59560
rect 3049 59530 3115 59533
rect 0 59528 3115 59530
rect 0 59472 3054 59528
rect 3110 59472 3115 59528
rect 0 59470 3115 59472
rect 0 59440 800 59470
rect 3049 59467 3115 59470
rect 10133 59530 10199 59533
rect 11200 59530 12000 59560
rect 10133 59528 12000 59530
rect 10133 59472 10138 59528
rect 10194 59472 12000 59528
rect 10133 59470 12000 59472
rect 10133 59467 10199 59470
rect 11200 59440 12000 59470
rect 2576 59328 2896 59329
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5839 59328 6159 59329
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 59263 6159 59264
rect 9103 59328 9423 59329
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 59263 9423 59264
rect 0 59122 800 59152
rect 1393 59122 1459 59125
rect 0 59120 1459 59122
rect 0 59064 1398 59120
rect 1454 59064 1459 59120
rect 0 59062 1459 59064
rect 0 59032 800 59062
rect 1393 59059 1459 59062
rect 1577 58850 1643 58853
rect 1894 58850 1900 58852
rect 1577 58848 1900 58850
rect 1577 58792 1582 58848
rect 1638 58792 1900 58848
rect 1577 58790 1900 58792
rect 1577 58787 1643 58790
rect 1894 58788 1900 58790
rect 1964 58788 1970 58852
rect 4207 58784 4527 58785
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 58719 4527 58720
rect 7471 58784 7791 58785
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 58719 7791 58720
rect 10133 58714 10199 58717
rect 11200 58714 12000 58744
rect 10133 58712 12000 58714
rect 10133 58656 10138 58712
rect 10194 58656 12000 58712
rect 10133 58654 12000 58656
rect 10133 58651 10199 58654
rect 11200 58624 12000 58654
rect 0 58578 800 58608
rect 1485 58578 1551 58581
rect 0 58576 1551 58578
rect 0 58520 1490 58576
rect 1546 58520 1551 58576
rect 0 58518 1551 58520
rect 0 58488 800 58518
rect 1485 58515 1551 58518
rect 1669 58578 1735 58581
rect 2313 58578 2379 58581
rect 1669 58576 2379 58578
rect 1669 58520 1674 58576
rect 1730 58520 2318 58576
rect 2374 58520 2379 58576
rect 1669 58518 2379 58520
rect 1669 58515 1735 58518
rect 2313 58515 2379 58518
rect 2576 58240 2896 58241
rect 0 58170 800 58200
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5839 58240 6159 58241
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 58175 6159 58176
rect 9103 58240 9423 58241
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 58175 9423 58176
rect 2405 58170 2471 58173
rect 0 58168 2471 58170
rect 0 58112 2410 58168
rect 2466 58112 2471 58168
rect 0 58110 2471 58112
rect 0 58080 800 58110
rect 2405 58107 2471 58110
rect 10133 58034 10199 58037
rect 11200 58034 12000 58064
rect 10133 58032 12000 58034
rect 10133 57976 10138 58032
rect 10194 57976 12000 58032
rect 10133 57974 12000 57976
rect 10133 57971 10199 57974
rect 11200 57944 12000 57974
rect 3049 57898 3115 57901
rect 3182 57898 3188 57900
rect 3049 57896 3188 57898
rect 3049 57840 3054 57896
rect 3110 57840 3188 57896
rect 3049 57838 3188 57840
rect 3049 57835 3115 57838
rect 3182 57836 3188 57838
rect 3252 57836 3258 57900
rect 0 57762 800 57792
rect 2773 57762 2839 57765
rect 0 57760 2839 57762
rect 0 57704 2778 57760
rect 2834 57704 2839 57760
rect 0 57702 2839 57704
rect 0 57672 800 57702
rect 2773 57699 2839 57702
rect 4207 57696 4527 57697
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 57631 4527 57632
rect 7471 57696 7791 57697
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 57631 7791 57632
rect 0 57354 800 57384
rect 2221 57354 2287 57357
rect 0 57352 2287 57354
rect 0 57296 2226 57352
rect 2282 57296 2287 57352
rect 0 57294 2287 57296
rect 0 57264 800 57294
rect 2221 57291 2287 57294
rect 10133 57218 10199 57221
rect 11200 57218 12000 57248
rect 10133 57216 12000 57218
rect 10133 57160 10138 57216
rect 10194 57160 12000 57216
rect 10133 57158 12000 57160
rect 10133 57155 10199 57158
rect 2576 57152 2896 57153
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5839 57152 6159 57153
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 57087 6159 57088
rect 9103 57152 9423 57153
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 11200 57128 12000 57158
rect 9103 57087 9423 57088
rect 0 56946 800 56976
rect 1485 56946 1551 56949
rect 0 56944 1551 56946
rect 0 56888 1490 56944
rect 1546 56888 1551 56944
rect 0 56886 1551 56888
rect 0 56856 800 56886
rect 1485 56883 1551 56886
rect 3366 56884 3372 56948
rect 3436 56946 3442 56948
rect 3509 56946 3575 56949
rect 3436 56944 3575 56946
rect 3436 56888 3514 56944
rect 3570 56888 3575 56944
rect 3436 56886 3575 56888
rect 3436 56884 3442 56886
rect 3509 56883 3575 56886
rect 4207 56608 4527 56609
rect 0 56538 800 56568
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 56543 4527 56544
rect 7471 56608 7791 56609
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 56543 7791 56544
rect 1485 56538 1551 56541
rect 0 56536 1551 56538
rect 0 56480 1490 56536
rect 1546 56480 1551 56536
rect 0 56478 1551 56480
rect 0 56448 800 56478
rect 1485 56475 1551 56478
rect 10133 56402 10199 56405
rect 11200 56402 12000 56432
rect 10133 56400 12000 56402
rect 10133 56344 10138 56400
rect 10194 56344 12000 56400
rect 10133 56342 12000 56344
rect 10133 56339 10199 56342
rect 11200 56312 12000 56342
rect 2576 56064 2896 56065
rect 0 55994 800 56024
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5839 56064 6159 56065
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 55999 6159 56000
rect 9103 56064 9423 56065
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 55999 9423 56000
rect 2221 55994 2287 55997
rect 0 55992 2287 55994
rect 0 55936 2226 55992
rect 2282 55936 2287 55992
rect 0 55934 2287 55936
rect 0 55904 800 55934
rect 2221 55931 2287 55934
rect 10133 55722 10199 55725
rect 11200 55722 12000 55752
rect 10133 55720 12000 55722
rect 10133 55664 10138 55720
rect 10194 55664 12000 55720
rect 10133 55662 12000 55664
rect 10133 55659 10199 55662
rect 11200 55632 12000 55662
rect 0 55586 800 55616
rect 2313 55586 2379 55589
rect 0 55584 2379 55586
rect 0 55528 2318 55584
rect 2374 55528 2379 55584
rect 0 55526 2379 55528
rect 0 55496 800 55526
rect 2313 55523 2379 55526
rect 4207 55520 4527 55521
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 55455 4527 55456
rect 7471 55520 7791 55521
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 55455 7791 55456
rect 1485 55450 1551 55453
rect 1485 55448 1594 55450
rect 1485 55392 1490 55448
rect 1546 55392 1594 55448
rect 1485 55387 1594 55392
rect 1393 55312 1459 55317
rect 1393 55256 1398 55312
rect 1454 55256 1459 55312
rect 1393 55251 1459 55256
rect 0 55178 800 55208
rect 1396 55178 1456 55251
rect 0 55118 1456 55178
rect 0 55088 800 55118
rect 0 54770 800 54800
rect 1534 54770 1594 55387
rect 2576 54976 2896 54977
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 5839 54976 6159 54977
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 54911 6159 54912
rect 9103 54976 9423 54977
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 54911 9423 54912
rect 10225 54906 10291 54909
rect 11200 54906 12000 54936
rect 10225 54904 12000 54906
rect 10225 54848 10230 54904
rect 10286 54848 12000 54904
rect 10225 54846 12000 54848
rect 10225 54843 10291 54846
rect 11200 54816 12000 54846
rect 0 54710 1594 54770
rect 0 54680 800 54710
rect 4207 54432 4527 54433
rect 0 54362 800 54392
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 54367 4527 54368
rect 7471 54432 7791 54433
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 54367 7791 54368
rect 2773 54362 2839 54365
rect 0 54360 2839 54362
rect 0 54304 2778 54360
rect 2834 54304 2839 54360
rect 0 54302 2839 54304
rect 0 54272 800 54302
rect 2773 54299 2839 54302
rect 10041 54090 10107 54093
rect 11200 54090 12000 54120
rect 10041 54088 12000 54090
rect 10041 54032 10046 54088
rect 10102 54032 12000 54088
rect 10041 54030 12000 54032
rect 10041 54027 10107 54030
rect 11200 54000 12000 54030
rect 0 53954 800 53984
rect 1393 53954 1459 53957
rect 0 53952 1459 53954
rect 0 53896 1398 53952
rect 1454 53896 1459 53952
rect 0 53894 1459 53896
rect 0 53864 800 53894
rect 1393 53891 1459 53894
rect 2576 53888 2896 53889
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5839 53888 6159 53889
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 53823 6159 53824
rect 9103 53888 9423 53889
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 53823 9423 53824
rect 0 53546 800 53576
rect 1485 53546 1551 53549
rect 0 53544 1551 53546
rect 0 53488 1490 53544
rect 1546 53488 1551 53544
rect 0 53486 1551 53488
rect 0 53456 800 53486
rect 1485 53483 1551 53486
rect 10041 53410 10107 53413
rect 11200 53410 12000 53440
rect 10041 53408 12000 53410
rect 10041 53352 10046 53408
rect 10102 53352 12000 53408
rect 10041 53350 12000 53352
rect 10041 53347 10107 53350
rect 4207 53344 4527 53345
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 53279 4527 53280
rect 7471 53344 7791 53345
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 11200 53320 12000 53350
rect 7471 53279 7791 53280
rect 0 53002 800 53032
rect 3049 53002 3115 53005
rect 0 53000 3115 53002
rect 0 52944 3054 53000
rect 3110 52944 3115 53000
rect 0 52942 3115 52944
rect 0 52912 800 52942
rect 3049 52939 3115 52942
rect 2576 52800 2896 52801
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 5839 52800 6159 52801
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 52735 6159 52736
rect 9103 52800 9423 52801
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 52735 9423 52736
rect 0 52594 800 52624
rect 2313 52594 2379 52597
rect 0 52592 2379 52594
rect 0 52536 2318 52592
rect 2374 52536 2379 52592
rect 0 52534 2379 52536
rect 0 52504 800 52534
rect 2313 52531 2379 52534
rect 10041 52594 10107 52597
rect 11200 52594 12000 52624
rect 10041 52592 12000 52594
rect 10041 52536 10046 52592
rect 10102 52536 12000 52592
rect 10041 52534 12000 52536
rect 10041 52531 10107 52534
rect 11200 52504 12000 52534
rect 4207 52256 4527 52257
rect 0 52186 800 52216
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 52191 4527 52192
rect 7471 52256 7791 52257
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 52191 7791 52192
rect 1393 52186 1459 52189
rect 0 52184 1459 52186
rect 0 52128 1398 52184
rect 1454 52128 1459 52184
rect 0 52126 1459 52128
rect 0 52096 800 52126
rect 1393 52123 1459 52126
rect 1669 51916 1735 51917
rect 1669 51914 1716 51916
rect 1624 51912 1716 51914
rect 1624 51856 1674 51912
rect 1624 51854 1716 51856
rect 1669 51852 1716 51854
rect 1780 51852 1786 51916
rect 1669 51851 1735 51852
rect 0 51778 800 51808
rect 1485 51778 1551 51781
rect 0 51776 1551 51778
rect 0 51720 1490 51776
rect 1546 51720 1551 51776
rect 0 51718 1551 51720
rect 0 51688 800 51718
rect 1485 51715 1551 51718
rect 10041 51778 10107 51781
rect 11200 51778 12000 51808
rect 10041 51776 12000 51778
rect 10041 51720 10046 51776
rect 10102 51720 12000 51776
rect 10041 51718 12000 51720
rect 10041 51715 10107 51718
rect 2576 51712 2896 51713
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 5839 51712 6159 51713
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 51647 6159 51648
rect 9103 51712 9423 51713
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 11200 51688 12000 51718
rect 9103 51647 9423 51648
rect 0 51370 800 51400
rect 3049 51370 3115 51373
rect 0 51368 3115 51370
rect 0 51312 3054 51368
rect 3110 51312 3115 51368
rect 0 51310 3115 51312
rect 0 51280 800 51310
rect 3049 51307 3115 51310
rect 4207 51168 4527 51169
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 51103 4527 51104
rect 7471 51168 7791 51169
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 51103 7791 51104
rect 10041 51098 10107 51101
rect 11200 51098 12000 51128
rect 10041 51096 12000 51098
rect 10041 51040 10046 51096
rect 10102 51040 12000 51096
rect 10041 51038 12000 51040
rect 10041 51035 10107 51038
rect 11200 51008 12000 51038
rect 0 50962 800 50992
rect 2221 50962 2287 50965
rect 0 50960 2287 50962
rect 0 50904 2226 50960
rect 2282 50904 2287 50960
rect 0 50902 2287 50904
rect 0 50872 800 50902
rect 2221 50899 2287 50902
rect 2576 50624 2896 50625
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 5839 50624 6159 50625
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 50559 6159 50560
rect 9103 50624 9423 50625
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 50559 9423 50560
rect 0 50418 800 50448
rect 1393 50418 1459 50421
rect 0 50416 1459 50418
rect 0 50360 1398 50416
rect 1454 50360 1459 50416
rect 0 50358 1459 50360
rect 0 50328 800 50358
rect 1393 50355 1459 50358
rect 3182 50356 3188 50420
rect 3252 50418 3258 50420
rect 3693 50418 3759 50421
rect 3252 50416 3759 50418
rect 3252 50360 3698 50416
rect 3754 50360 3759 50416
rect 3252 50358 3759 50360
rect 3252 50356 3258 50358
rect 3693 50355 3759 50358
rect 4613 50420 4679 50421
rect 4613 50416 4660 50420
rect 4724 50418 4730 50420
rect 4613 50360 4618 50416
rect 4613 50356 4660 50360
rect 4724 50358 4770 50418
rect 4724 50356 4730 50358
rect 4613 50355 4679 50356
rect 10041 50282 10107 50285
rect 11200 50282 12000 50312
rect 10041 50280 12000 50282
rect 10041 50224 10046 50280
rect 10102 50224 12000 50280
rect 10041 50222 12000 50224
rect 10041 50219 10107 50222
rect 11200 50192 12000 50222
rect 4207 50080 4527 50081
rect 0 50010 800 50040
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 50015 4527 50016
rect 7471 50080 7791 50081
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 50015 7791 50016
rect 1485 50010 1551 50013
rect 0 50008 1551 50010
rect 0 49952 1490 50008
rect 1546 49952 1551 50008
rect 0 49950 1551 49952
rect 0 49920 800 49950
rect 1485 49947 1551 49950
rect 0 49602 800 49632
rect 2405 49602 2471 49605
rect 0 49600 2471 49602
rect 0 49544 2410 49600
rect 2466 49544 2471 49600
rect 0 49542 2471 49544
rect 0 49512 800 49542
rect 2405 49539 2471 49542
rect 2576 49536 2896 49537
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 5839 49536 6159 49537
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 49471 6159 49472
rect 9103 49536 9423 49537
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 49471 9423 49472
rect 10041 49466 10107 49469
rect 11200 49466 12000 49496
rect 10041 49464 12000 49466
rect 10041 49408 10046 49464
rect 10102 49408 12000 49464
rect 10041 49406 12000 49408
rect 10041 49403 10107 49406
rect 11200 49376 12000 49406
rect 0 49194 800 49224
rect 2221 49194 2287 49197
rect 0 49192 2287 49194
rect 0 49136 2226 49192
rect 2282 49136 2287 49192
rect 0 49134 2287 49136
rect 0 49104 800 49134
rect 2221 49131 2287 49134
rect 4207 48992 4527 48993
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 48927 4527 48928
rect 7471 48992 7791 48993
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 48927 7791 48928
rect 0 48786 800 48816
rect 2773 48786 2839 48789
rect 0 48784 2839 48786
rect 0 48728 2778 48784
rect 2834 48728 2839 48784
rect 0 48726 2839 48728
rect 0 48696 800 48726
rect 2773 48723 2839 48726
rect 4521 48786 4587 48789
rect 4654 48786 4660 48788
rect 4521 48784 4660 48786
rect 4521 48728 4526 48784
rect 4582 48728 4660 48784
rect 4521 48726 4660 48728
rect 4521 48723 4587 48726
rect 4654 48724 4660 48726
rect 4724 48724 4730 48788
rect 10041 48786 10107 48789
rect 11200 48786 12000 48816
rect 10041 48784 12000 48786
rect 10041 48728 10046 48784
rect 10102 48728 12000 48784
rect 10041 48726 12000 48728
rect 10041 48723 10107 48726
rect 11200 48696 12000 48726
rect 2576 48448 2896 48449
rect 0 48378 800 48408
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 5839 48448 6159 48449
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 48383 6159 48384
rect 9103 48448 9423 48449
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 48383 9423 48384
rect 1485 48378 1551 48381
rect 1945 48380 2011 48381
rect 1894 48378 1900 48380
rect 0 48376 1551 48378
rect 0 48320 1490 48376
rect 1546 48320 1551 48376
rect 0 48318 1551 48320
rect 1854 48318 1900 48378
rect 1964 48376 2011 48380
rect 3366 48378 3372 48380
rect 2006 48320 2011 48376
rect 3006 48333 3372 48378
rect 0 48288 800 48318
rect 1485 48315 1551 48318
rect 1894 48316 1900 48318
rect 1964 48316 2011 48320
rect 1945 48315 2011 48316
rect 2957 48328 3372 48333
rect 2957 48272 2962 48328
rect 3018 48318 3372 48328
rect 3018 48272 3066 48318
rect 3366 48316 3372 48318
rect 3436 48316 3442 48380
rect 2957 48270 3066 48272
rect 2957 48267 3023 48270
rect 10041 47970 10107 47973
rect 11200 47970 12000 48000
rect 10041 47968 12000 47970
rect 10041 47912 10046 47968
rect 10102 47912 12000 47968
rect 10041 47910 12000 47912
rect 10041 47907 10107 47910
rect 4207 47904 4527 47905
rect 0 47834 800 47864
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 47839 4527 47840
rect 7471 47904 7791 47905
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 11200 47880 12000 47910
rect 7471 47839 7791 47840
rect 1485 47834 1551 47837
rect 0 47832 1551 47834
rect 0 47776 1490 47832
rect 1546 47776 1551 47832
rect 0 47774 1551 47776
rect 0 47744 800 47774
rect 1485 47771 1551 47774
rect 2773 47834 2839 47837
rect 2998 47834 3004 47836
rect 2773 47832 3004 47834
rect 2773 47776 2778 47832
rect 2834 47776 3004 47832
rect 2773 47774 3004 47776
rect 2773 47771 2839 47774
rect 2998 47772 3004 47774
rect 3068 47834 3074 47836
rect 3509 47834 3575 47837
rect 3068 47832 3575 47834
rect 3068 47776 3514 47832
rect 3570 47776 3575 47832
rect 3068 47774 3575 47776
rect 3068 47772 3074 47774
rect 3509 47771 3575 47774
rect 1485 47562 1551 47565
rect 1166 47560 1551 47562
rect 1166 47504 1490 47560
rect 1546 47504 1551 47560
rect 1166 47502 1551 47504
rect 0 47426 800 47456
rect 1166 47426 1226 47502
rect 1485 47499 1551 47502
rect 2681 47562 2747 47565
rect 4654 47562 4660 47564
rect 2681 47560 4660 47562
rect 2681 47504 2686 47560
rect 2742 47504 4660 47560
rect 2681 47502 4660 47504
rect 2681 47499 2747 47502
rect 4654 47500 4660 47502
rect 4724 47500 4730 47564
rect 5901 47562 5967 47565
rect 6310 47562 6316 47564
rect 5901 47560 6316 47562
rect 5901 47504 5906 47560
rect 5962 47504 6316 47560
rect 5901 47502 6316 47504
rect 5901 47499 5967 47502
rect 6310 47500 6316 47502
rect 6380 47500 6386 47564
rect 0 47366 1226 47426
rect 0 47336 800 47366
rect 2576 47360 2896 47361
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 5839 47360 6159 47361
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 47295 6159 47296
rect 9103 47360 9423 47361
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 47295 9423 47296
rect 2078 47092 2084 47156
rect 2148 47154 2154 47156
rect 3693 47154 3759 47157
rect 2148 47152 3759 47154
rect 2148 47096 3698 47152
rect 3754 47096 3759 47152
rect 2148 47094 3759 47096
rect 2148 47092 2154 47094
rect 3693 47091 3759 47094
rect 10041 47154 10107 47157
rect 11200 47154 12000 47184
rect 10041 47152 12000 47154
rect 10041 47096 10046 47152
rect 10102 47096 12000 47152
rect 10041 47094 12000 47096
rect 10041 47091 10107 47094
rect 11200 47064 12000 47094
rect 0 47018 800 47048
rect 1485 47018 1551 47021
rect 0 47016 1551 47018
rect 0 46960 1490 47016
rect 1546 46960 1551 47016
rect 0 46958 1551 46960
rect 0 46928 800 46958
rect 1485 46955 1551 46958
rect 4207 46816 4527 46817
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 46751 4527 46752
rect 7471 46816 7791 46817
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 46751 7791 46752
rect 0 46610 800 46640
rect 1485 46610 1551 46613
rect 0 46608 1551 46610
rect 0 46552 1490 46608
rect 1546 46552 1551 46608
rect 0 46550 1551 46552
rect 0 46520 800 46550
rect 1485 46547 1551 46550
rect 2773 46474 2839 46477
rect 2998 46474 3004 46476
rect 2773 46472 3004 46474
rect 2773 46416 2778 46472
rect 2834 46416 3004 46472
rect 2773 46414 3004 46416
rect 2773 46411 2839 46414
rect 2998 46412 3004 46414
rect 3068 46412 3074 46476
rect 10041 46474 10107 46477
rect 11200 46474 12000 46504
rect 10041 46472 12000 46474
rect 10041 46416 10046 46472
rect 10102 46416 12000 46472
rect 10041 46414 12000 46416
rect 10041 46411 10107 46414
rect 11200 46384 12000 46414
rect 2576 46272 2896 46273
rect 0 46202 800 46232
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 5839 46272 6159 46273
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 46207 6159 46208
rect 9103 46272 9423 46273
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 46207 9423 46208
rect 1485 46202 1551 46205
rect 0 46200 1551 46202
rect 0 46144 1490 46200
rect 1546 46144 1551 46200
rect 0 46142 1551 46144
rect 0 46112 800 46142
rect 1485 46139 1551 46142
rect 4429 46066 4495 46069
rect 4429 46064 5090 46066
rect 4429 46008 4434 46064
rect 4490 46008 5090 46064
rect 4429 46006 5090 46008
rect 4429 46003 4495 46006
rect 1577 45930 1643 45933
rect 1577 45928 1778 45930
rect 1577 45872 1582 45928
rect 1638 45872 1778 45928
rect 1577 45870 1778 45872
rect 1577 45867 1643 45870
rect 0 45794 800 45824
rect 1485 45794 1551 45797
rect 0 45792 1551 45794
rect 0 45736 1490 45792
rect 1546 45736 1551 45792
rect 0 45734 1551 45736
rect 0 45704 800 45734
rect 1485 45731 1551 45734
rect 0 45250 800 45280
rect 0 45190 1410 45250
rect 0 45160 800 45190
rect 1350 44978 1410 45190
rect 1718 45114 1778 45870
rect 4207 45728 4527 45729
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 45663 4527 45664
rect 5030 45522 5090 46006
rect 7471 45728 7791 45729
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 45663 7791 45664
rect 10041 45658 10107 45661
rect 11200 45658 12000 45688
rect 10041 45656 12000 45658
rect 10041 45600 10046 45656
rect 10102 45600 12000 45656
rect 10041 45598 12000 45600
rect 10041 45595 10107 45598
rect 11200 45568 12000 45598
rect 5165 45522 5231 45525
rect 5030 45520 5231 45522
rect 5030 45464 5170 45520
rect 5226 45464 5231 45520
rect 5030 45462 5231 45464
rect 5165 45459 5231 45462
rect 2221 45386 2287 45389
rect 3417 45386 3483 45389
rect 2221 45384 3483 45386
rect 2221 45328 2226 45384
rect 2282 45328 3422 45384
rect 3478 45328 3483 45384
rect 2221 45326 3483 45328
rect 2221 45323 2287 45326
rect 3417 45323 3483 45326
rect 2576 45184 2896 45185
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 5839 45184 6159 45185
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 45119 6159 45120
rect 9103 45184 9423 45185
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 45119 9423 45120
rect 1853 45114 1919 45117
rect 1718 45112 1919 45114
rect 1718 45056 1858 45112
rect 1914 45056 1919 45112
rect 1718 45054 1919 45056
rect 1853 45051 1919 45054
rect 2773 44978 2839 44981
rect 1350 44976 2839 44978
rect 1350 44920 2778 44976
rect 2834 44920 2839 44976
rect 1350 44918 2839 44920
rect 2773 44915 2839 44918
rect 0 44842 800 44872
rect 1485 44842 1551 44845
rect 0 44840 1551 44842
rect 0 44784 1490 44840
rect 1546 44784 1551 44840
rect 0 44782 1551 44784
rect 0 44752 800 44782
rect 1485 44779 1551 44782
rect 10041 44842 10107 44845
rect 11200 44842 12000 44872
rect 10041 44840 12000 44842
rect 10041 44784 10046 44840
rect 10102 44784 12000 44840
rect 10041 44782 12000 44784
rect 10041 44779 10107 44782
rect 11200 44752 12000 44782
rect 4207 44640 4527 44641
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 44575 4527 44576
rect 7471 44640 7791 44641
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 44575 7791 44576
rect 0 44434 800 44464
rect 2773 44434 2839 44437
rect 0 44432 2839 44434
rect 0 44376 2778 44432
rect 2834 44376 2839 44432
rect 0 44374 2839 44376
rect 0 44344 800 44374
rect 2773 44371 2839 44374
rect 2998 44372 3004 44436
rect 3068 44434 3074 44436
rect 4153 44434 4219 44437
rect 3068 44432 4219 44434
rect 3068 44376 4158 44432
rect 4214 44376 4219 44432
rect 3068 44374 4219 44376
rect 3068 44372 3074 44374
rect 4153 44371 4219 44374
rect 10041 44162 10107 44165
rect 11200 44162 12000 44192
rect 10041 44160 12000 44162
rect 10041 44104 10046 44160
rect 10102 44104 12000 44160
rect 10041 44102 12000 44104
rect 10041 44099 10107 44102
rect 2576 44096 2896 44097
rect 0 44026 800 44056
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5839 44096 6159 44097
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 44031 6159 44032
rect 9103 44096 9423 44097
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 11200 44072 12000 44102
rect 9103 44031 9423 44032
rect 0 43966 1410 44026
rect 0 43936 800 43966
rect 1350 43890 1410 43966
rect 2957 43890 3023 43893
rect 1350 43888 3023 43890
rect 1350 43832 2962 43888
rect 3018 43832 3023 43888
rect 1350 43830 3023 43832
rect 2957 43827 3023 43830
rect 6310 43692 6316 43756
rect 6380 43754 6386 43756
rect 6729 43754 6795 43757
rect 6380 43752 6795 43754
rect 6380 43696 6734 43752
rect 6790 43696 6795 43752
rect 6380 43694 6795 43696
rect 6380 43692 6386 43694
rect 6729 43691 6795 43694
rect 0 43618 800 43648
rect 2313 43618 2379 43621
rect 0 43616 2379 43618
rect 0 43560 2318 43616
rect 2374 43560 2379 43616
rect 0 43558 2379 43560
rect 0 43528 800 43558
rect 2313 43555 2379 43558
rect 4207 43552 4527 43553
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 43487 4527 43488
rect 7471 43552 7791 43553
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 43487 7791 43488
rect 10041 43346 10107 43349
rect 11200 43346 12000 43376
rect 10041 43344 12000 43346
rect 10041 43288 10046 43344
rect 10102 43288 12000 43344
rect 10041 43286 12000 43288
rect 10041 43283 10107 43286
rect 11200 43256 12000 43286
rect 0 43210 800 43240
rect 2773 43210 2839 43213
rect 0 43208 2839 43210
rect 0 43152 2778 43208
rect 2834 43152 2839 43208
rect 0 43150 2839 43152
rect 0 43120 800 43150
rect 2773 43147 2839 43150
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 5839 43008 6159 43009
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 42943 6159 42944
rect 9103 43008 9423 43009
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 42943 9423 42944
rect 0 42666 800 42696
rect 2957 42666 3023 42669
rect 0 42664 3023 42666
rect 0 42608 2962 42664
rect 3018 42608 3023 42664
rect 0 42606 3023 42608
rect 0 42576 800 42606
rect 2957 42603 3023 42606
rect 4654 42468 4660 42532
rect 4724 42530 4730 42532
rect 5073 42530 5139 42533
rect 4724 42528 5139 42530
rect 4724 42472 5078 42528
rect 5134 42472 5139 42528
rect 4724 42470 5139 42472
rect 4724 42468 4730 42470
rect 5073 42467 5139 42470
rect 10041 42530 10107 42533
rect 11200 42530 12000 42560
rect 10041 42528 12000 42530
rect 10041 42472 10046 42528
rect 10102 42472 12000 42528
rect 10041 42470 12000 42472
rect 10041 42467 10107 42470
rect 4207 42464 4527 42465
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 42399 4527 42400
rect 7471 42464 7791 42465
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 11200 42440 12000 42470
rect 7471 42399 7791 42400
rect 0 42258 800 42288
rect 3049 42258 3115 42261
rect 0 42256 3115 42258
rect 0 42200 3054 42256
rect 3110 42200 3115 42256
rect 0 42198 3115 42200
rect 0 42168 800 42198
rect 3049 42195 3115 42198
rect 2576 41920 2896 41921
rect 0 41850 800 41880
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5839 41920 6159 41921
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 41855 6159 41856
rect 9103 41920 9423 41921
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 41855 9423 41856
rect 2221 41850 2287 41853
rect 0 41848 2287 41850
rect 0 41792 2226 41848
rect 2282 41792 2287 41848
rect 0 41790 2287 41792
rect 0 41760 800 41790
rect 2221 41787 2287 41790
rect 10041 41850 10107 41853
rect 11200 41850 12000 41880
rect 10041 41848 12000 41850
rect 10041 41792 10046 41848
rect 10102 41792 12000 41848
rect 10041 41790 12000 41792
rect 10041 41787 10107 41790
rect 11200 41760 12000 41790
rect 2998 41516 3004 41580
rect 3068 41578 3074 41580
rect 3417 41578 3483 41581
rect 3068 41576 3483 41578
rect 3068 41520 3422 41576
rect 3478 41520 3483 41576
rect 3068 41518 3483 41520
rect 3068 41516 3074 41518
rect 3417 41515 3483 41518
rect 0 41442 800 41472
rect 1485 41442 1551 41445
rect 0 41440 1551 41442
rect 0 41384 1490 41440
rect 1546 41384 1551 41440
rect 0 41382 1551 41384
rect 0 41352 800 41382
rect 1485 41379 1551 41382
rect 3601 41442 3667 41445
rect 3969 41442 4035 41445
rect 3601 41440 4035 41442
rect 3601 41384 3606 41440
rect 3662 41384 3974 41440
rect 4030 41384 4035 41440
rect 3601 41382 4035 41384
rect 3601 41379 3667 41382
rect 3969 41379 4035 41382
rect 4207 41376 4527 41377
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 41311 4527 41312
rect 7471 41376 7791 41377
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 41311 7791 41312
rect 2262 41108 2268 41172
rect 2332 41170 2338 41172
rect 2589 41170 2655 41173
rect 2332 41168 2655 41170
rect 2332 41112 2594 41168
rect 2650 41112 2655 41168
rect 2332 41110 2655 41112
rect 2332 41108 2338 41110
rect 2589 41107 2655 41110
rect 2998 41108 3004 41172
rect 3068 41170 3074 41172
rect 3325 41170 3391 41173
rect 3068 41168 3391 41170
rect 3068 41112 3330 41168
rect 3386 41112 3391 41168
rect 3068 41110 3391 41112
rect 3068 41108 3074 41110
rect 3325 41107 3391 41110
rect 0 41034 800 41064
rect 3049 41034 3115 41037
rect 0 41032 3115 41034
rect 0 40976 3054 41032
rect 3110 40976 3115 41032
rect 0 40974 3115 40976
rect 0 40944 800 40974
rect 3049 40971 3115 40974
rect 10041 41034 10107 41037
rect 11200 41034 12000 41064
rect 10041 41032 12000 41034
rect 10041 40976 10046 41032
rect 10102 40976 12000 41032
rect 10041 40974 12000 40976
rect 10041 40971 10107 40974
rect 11200 40944 12000 40974
rect 1945 40898 2011 40901
rect 2078 40898 2084 40900
rect 1945 40896 2084 40898
rect 1945 40840 1950 40896
rect 2006 40840 2084 40896
rect 1945 40838 2084 40840
rect 1945 40835 2011 40838
rect 2078 40836 2084 40838
rect 2148 40836 2154 40900
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5839 40832 6159 40833
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 40767 6159 40768
rect 9103 40832 9423 40833
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 40767 9423 40768
rect 0 40626 800 40656
rect 2221 40626 2287 40629
rect 0 40624 2287 40626
rect 0 40568 2226 40624
rect 2282 40568 2287 40624
rect 0 40566 2287 40568
rect 0 40536 800 40566
rect 2221 40563 2287 40566
rect 10041 40354 10107 40357
rect 11200 40354 12000 40384
rect 10041 40352 12000 40354
rect 10041 40296 10046 40352
rect 10102 40296 12000 40352
rect 10041 40294 12000 40296
rect 10041 40291 10107 40294
rect 4207 40288 4527 40289
rect 0 40218 800 40248
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 40223 4527 40224
rect 7471 40288 7791 40289
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 11200 40264 12000 40294
rect 7471 40223 7791 40224
rect 1209 40218 1275 40221
rect 0 40216 1275 40218
rect 0 40160 1214 40216
rect 1270 40160 1275 40216
rect 0 40158 1275 40160
rect 0 40128 800 40158
rect 1209 40155 1275 40158
rect 1894 40020 1900 40084
rect 1964 40082 1970 40084
rect 2129 40082 2195 40085
rect 1964 40080 2195 40082
rect 1964 40024 2134 40080
rect 2190 40024 2195 40080
rect 1964 40022 2195 40024
rect 1964 40020 1970 40022
rect 2129 40019 2195 40022
rect 2576 39744 2896 39745
rect 0 39674 800 39704
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 5839 39744 6159 39745
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 39679 6159 39680
rect 9103 39744 9423 39745
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 39679 9423 39680
rect 1485 39674 1551 39677
rect 0 39672 1551 39674
rect 0 39616 1490 39672
rect 1546 39616 1551 39672
rect 0 39614 1551 39616
rect 0 39584 800 39614
rect 1485 39611 1551 39614
rect 10041 39538 10107 39541
rect 11200 39538 12000 39568
rect 10041 39536 12000 39538
rect 10041 39480 10046 39536
rect 10102 39480 12000 39536
rect 10041 39478 12000 39480
rect 10041 39475 10107 39478
rect 11200 39448 12000 39478
rect 0 39266 800 39296
rect 2773 39266 2839 39269
rect 0 39264 2839 39266
rect 0 39208 2778 39264
rect 2834 39208 2839 39264
rect 0 39206 2839 39208
rect 0 39176 800 39206
rect 2773 39203 2839 39206
rect 4207 39200 4527 39201
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 39135 4527 39136
rect 7471 39200 7791 39201
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 39135 7791 39136
rect 0 38858 800 38888
rect 1209 38858 1275 38861
rect 0 38856 1275 38858
rect 0 38800 1214 38856
rect 1270 38800 1275 38856
rect 0 38798 1275 38800
rect 0 38768 800 38798
rect 1209 38795 1275 38798
rect 10041 38722 10107 38725
rect 11200 38722 12000 38752
rect 10041 38720 12000 38722
rect 10041 38664 10046 38720
rect 10102 38664 12000 38720
rect 10041 38662 12000 38664
rect 10041 38659 10107 38662
rect 2576 38656 2896 38657
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 5839 38656 6159 38657
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 38591 6159 38592
rect 9103 38656 9423 38657
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 11200 38632 12000 38662
rect 9103 38591 9423 38592
rect 0 38450 800 38480
rect 3417 38450 3483 38453
rect 0 38448 3483 38450
rect 0 38392 3422 38448
rect 3478 38392 3483 38448
rect 0 38390 3483 38392
rect 0 38360 800 38390
rect 3417 38387 3483 38390
rect 3601 38314 3667 38317
rect 3734 38314 3740 38316
rect 3601 38312 3740 38314
rect 3601 38256 3606 38312
rect 3662 38256 3740 38312
rect 3601 38254 3740 38256
rect 3601 38251 3667 38254
rect 3734 38252 3740 38254
rect 3804 38252 3810 38316
rect 4207 38112 4527 38113
rect 0 38042 800 38072
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 38047 4527 38048
rect 7471 38112 7791 38113
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 38047 7791 38048
rect 2957 38042 3023 38045
rect 0 38040 3023 38042
rect 0 37984 2962 38040
rect 3018 37984 3023 38040
rect 0 37982 3023 37984
rect 0 37952 800 37982
rect 2957 37979 3023 37982
rect 10041 38042 10107 38045
rect 11200 38042 12000 38072
rect 10041 38040 12000 38042
rect 10041 37984 10046 38040
rect 10102 37984 12000 38040
rect 10041 37982 12000 37984
rect 10041 37979 10107 37982
rect 11200 37952 12000 37982
rect 1485 37768 1551 37773
rect 1485 37712 1490 37768
rect 1546 37712 1551 37768
rect 1485 37707 1551 37712
rect 0 37634 800 37664
rect 1488 37634 1548 37707
rect 0 37574 1548 37634
rect 0 37544 800 37574
rect 2576 37568 2896 37569
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5839 37568 6159 37569
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 37503 6159 37504
rect 9103 37568 9423 37569
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 37503 9423 37504
rect 3233 37362 3299 37365
rect 3366 37362 3372 37364
rect 3233 37360 3372 37362
rect 3233 37304 3238 37360
rect 3294 37304 3372 37360
rect 3233 37302 3372 37304
rect 3233 37299 3299 37302
rect 3366 37300 3372 37302
rect 3436 37300 3442 37364
rect 10041 37226 10107 37229
rect 11200 37226 12000 37256
rect 10041 37224 12000 37226
rect 10041 37168 10046 37224
rect 10102 37168 12000 37224
rect 10041 37166 12000 37168
rect 10041 37163 10107 37166
rect 11200 37136 12000 37166
rect 0 37090 800 37120
rect 1485 37090 1551 37093
rect 0 37088 1551 37090
rect 0 37032 1490 37088
rect 1546 37032 1551 37088
rect 0 37030 1551 37032
rect 0 37000 800 37030
rect 1485 37027 1551 37030
rect 2221 37090 2287 37093
rect 2221 37088 2330 37090
rect 2221 37032 2226 37088
rect 2282 37032 2330 37088
rect 2221 37027 2330 37032
rect 2270 36821 2330 37027
rect 4207 37024 4527 37025
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 36959 4527 36960
rect 7471 37024 7791 37025
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 36959 7791 36960
rect 2221 36816 2330 36821
rect 2221 36760 2226 36816
rect 2282 36760 2330 36816
rect 2221 36758 2330 36760
rect 2221 36755 2287 36758
rect 0 36682 800 36712
rect 3049 36682 3115 36685
rect 0 36680 3115 36682
rect 0 36624 3054 36680
rect 3110 36624 3115 36680
rect 0 36622 3115 36624
rect 0 36592 800 36622
rect 3049 36619 3115 36622
rect 2576 36480 2896 36481
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 5839 36480 6159 36481
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 36415 6159 36416
rect 9103 36480 9423 36481
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 36415 9423 36416
rect 10041 36410 10107 36413
rect 11200 36410 12000 36440
rect 10041 36408 12000 36410
rect 10041 36352 10046 36408
rect 10102 36352 12000 36408
rect 10041 36350 12000 36352
rect 10041 36347 10107 36350
rect 11200 36320 12000 36350
rect 0 36274 800 36304
rect 2313 36274 2379 36277
rect 0 36272 2379 36274
rect 0 36216 2318 36272
rect 2374 36216 2379 36272
rect 0 36214 2379 36216
rect 0 36184 800 36214
rect 2313 36211 2379 36214
rect 4207 35936 4527 35937
rect 0 35866 800 35896
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 35871 4527 35872
rect 7471 35936 7791 35937
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 35871 7791 35872
rect 1485 35866 1551 35869
rect 0 35864 1551 35866
rect 0 35808 1490 35864
rect 1546 35808 1551 35864
rect 0 35806 1551 35808
rect 0 35776 800 35806
rect 1485 35803 1551 35806
rect 10041 35730 10107 35733
rect 11200 35730 12000 35760
rect 10041 35728 12000 35730
rect 10041 35672 10046 35728
rect 10102 35672 12000 35728
rect 10041 35670 12000 35672
rect 10041 35667 10107 35670
rect 11200 35640 12000 35670
rect 3049 35594 3115 35597
rect 1350 35592 3115 35594
rect 1350 35536 3054 35592
rect 3110 35536 3115 35592
rect 1350 35534 3115 35536
rect 0 35458 800 35488
rect 1350 35458 1410 35534
rect 3049 35531 3115 35534
rect 0 35398 1410 35458
rect 0 35368 800 35398
rect 2576 35392 2896 35393
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5839 35392 6159 35393
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 35327 6159 35328
rect 9103 35392 9423 35393
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 35327 9423 35328
rect 0 35050 800 35080
rect 1485 35050 1551 35053
rect 0 35048 1551 35050
rect 0 34992 1490 35048
rect 1546 34992 1551 35048
rect 0 34990 1551 34992
rect 0 34960 800 34990
rect 1485 34987 1551 34990
rect 10041 34914 10107 34917
rect 11200 34914 12000 34944
rect 10041 34912 12000 34914
rect 10041 34856 10046 34912
rect 10102 34856 12000 34912
rect 10041 34854 12000 34856
rect 10041 34851 10107 34854
rect 4207 34848 4527 34849
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 34783 4527 34784
rect 7471 34848 7791 34849
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 11200 34824 12000 34854
rect 7471 34783 7791 34784
rect 0 34506 800 34536
rect 3233 34506 3299 34509
rect 0 34504 3299 34506
rect 0 34448 3238 34504
rect 3294 34448 3299 34504
rect 0 34446 3299 34448
rect 0 34416 800 34446
rect 3233 34443 3299 34446
rect 2576 34304 2896 34305
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5839 34304 6159 34305
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 34239 6159 34240
rect 9103 34304 9423 34305
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 34239 9423 34240
rect 0 34098 800 34128
rect 2405 34098 2471 34101
rect 0 34096 2471 34098
rect 0 34040 2410 34096
rect 2466 34040 2471 34096
rect 0 34038 2471 34040
rect 0 34008 800 34038
rect 2405 34035 2471 34038
rect 10041 34098 10107 34101
rect 11200 34098 12000 34128
rect 10041 34096 12000 34098
rect 10041 34040 10046 34096
rect 10102 34040 12000 34096
rect 10041 34038 12000 34040
rect 10041 34035 10107 34038
rect 11200 34008 12000 34038
rect 4207 33760 4527 33761
rect 0 33690 800 33720
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 33695 4527 33696
rect 7471 33760 7791 33761
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 33695 7791 33696
rect 2313 33690 2379 33693
rect 0 33688 2379 33690
rect 0 33632 2318 33688
rect 2374 33632 2379 33688
rect 0 33630 2379 33632
rect 0 33600 800 33630
rect 2313 33627 2379 33630
rect 3366 33492 3372 33556
rect 3436 33554 3442 33556
rect 3509 33554 3575 33557
rect 3436 33552 3575 33554
rect 3436 33496 3514 33552
rect 3570 33496 3575 33552
rect 3436 33494 3575 33496
rect 3436 33492 3442 33494
rect 3509 33491 3575 33494
rect 10041 33418 10107 33421
rect 11200 33418 12000 33448
rect 10041 33416 12000 33418
rect 10041 33360 10046 33416
rect 10102 33360 12000 33416
rect 10041 33358 12000 33360
rect 10041 33355 10107 33358
rect 11200 33328 12000 33358
rect 0 33282 800 33312
rect 2313 33282 2379 33285
rect 0 33280 2379 33282
rect 0 33224 2318 33280
rect 2374 33224 2379 33280
rect 0 33222 2379 33224
rect 0 33192 800 33222
rect 2313 33219 2379 33222
rect 2576 33216 2896 33217
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5839 33216 6159 33217
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 33151 6159 33152
rect 9103 33216 9423 33217
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 33151 9423 33152
rect 0 32874 800 32904
rect 2313 32874 2379 32877
rect 0 32872 2379 32874
rect 0 32816 2318 32872
rect 2374 32816 2379 32872
rect 0 32814 2379 32816
rect 0 32784 800 32814
rect 2313 32811 2379 32814
rect 4207 32672 4527 32673
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 32607 4527 32608
rect 7471 32672 7791 32673
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 32607 7791 32608
rect 10041 32602 10107 32605
rect 11200 32602 12000 32632
rect 10041 32600 12000 32602
rect 10041 32544 10046 32600
rect 10102 32544 12000 32600
rect 10041 32542 12000 32544
rect 10041 32539 10107 32542
rect 11200 32512 12000 32542
rect 0 32466 800 32496
rect 1485 32466 1551 32469
rect 0 32464 1551 32466
rect 0 32408 1490 32464
rect 1546 32408 1551 32464
rect 0 32406 1551 32408
rect 0 32376 800 32406
rect 1485 32403 1551 32406
rect 2576 32128 2896 32129
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 5839 32128 6159 32129
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 32063 6159 32064
rect 9103 32128 9423 32129
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 32063 9423 32064
rect 2998 31996 3004 32060
rect 3068 32058 3074 32060
rect 3785 32058 3851 32061
rect 3068 32056 3851 32058
rect 3068 32000 3790 32056
rect 3846 32000 3851 32056
rect 3068 31998 3851 32000
rect 3068 31996 3074 31998
rect 3785 31995 3851 31998
rect 0 31922 800 31952
rect 1577 31922 1643 31925
rect 0 31920 1643 31922
rect 0 31864 1582 31920
rect 1638 31864 1643 31920
rect 0 31862 1643 31864
rect 0 31832 800 31862
rect 1577 31859 1643 31862
rect 1853 31924 1919 31925
rect 1853 31920 1900 31924
rect 1964 31922 1970 31924
rect 1853 31864 1858 31920
rect 1853 31860 1900 31864
rect 1964 31862 2010 31922
rect 1964 31860 1970 31862
rect 1853 31859 1919 31860
rect 1853 31786 1919 31789
rect 2262 31786 2268 31788
rect 1853 31784 2268 31786
rect 1853 31728 1858 31784
rect 1914 31728 2268 31784
rect 1853 31726 2268 31728
rect 1853 31723 1919 31726
rect 2262 31724 2268 31726
rect 2332 31724 2338 31788
rect 10041 31786 10107 31789
rect 11200 31786 12000 31816
rect 10041 31784 12000 31786
rect 10041 31728 10046 31784
rect 10102 31728 12000 31784
rect 10041 31726 12000 31728
rect 10041 31723 10107 31726
rect 11200 31696 12000 31726
rect 4207 31584 4527 31585
rect 0 31514 800 31544
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 31519 4527 31520
rect 7471 31584 7791 31585
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 31519 7791 31520
rect 2773 31514 2839 31517
rect 0 31512 2839 31514
rect 0 31456 2778 31512
rect 2834 31456 2839 31512
rect 0 31454 2839 31456
rect 0 31424 800 31454
rect 2773 31451 2839 31454
rect 0 31106 800 31136
rect 1485 31106 1551 31109
rect 0 31104 1551 31106
rect 0 31048 1490 31104
rect 1546 31048 1551 31104
rect 0 31046 1551 31048
rect 0 31016 800 31046
rect 1485 31043 1551 31046
rect 10041 31106 10107 31109
rect 11200 31106 12000 31136
rect 10041 31104 12000 31106
rect 10041 31048 10046 31104
rect 10102 31048 12000 31104
rect 10041 31046 12000 31048
rect 10041 31043 10107 31046
rect 2576 31040 2896 31041
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5839 31040 6159 31041
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 30975 6159 30976
rect 9103 31040 9423 31041
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 11200 31016 12000 31046
rect 9103 30975 9423 30976
rect 0 30698 800 30728
rect 1485 30698 1551 30701
rect 0 30696 1551 30698
rect 0 30640 1490 30696
rect 1546 30640 1551 30696
rect 0 30638 1551 30640
rect 0 30608 800 30638
rect 1485 30635 1551 30638
rect 4207 30496 4527 30497
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 30431 4527 30432
rect 7471 30496 7791 30497
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 30431 7791 30432
rect 0 30290 800 30320
rect 3969 30290 4035 30293
rect 0 30288 4035 30290
rect 0 30232 3974 30288
rect 4030 30232 4035 30288
rect 0 30230 4035 30232
rect 0 30200 800 30230
rect 3969 30227 4035 30230
rect 10041 30290 10107 30293
rect 11200 30290 12000 30320
rect 10041 30288 12000 30290
rect 10041 30232 10046 30288
rect 10102 30232 12000 30288
rect 10041 30230 12000 30232
rect 10041 30227 10107 30230
rect 11200 30200 12000 30230
rect 3785 30156 3851 30157
rect 3734 30154 3740 30156
rect 3694 30094 3740 30154
rect 3804 30152 3851 30156
rect 3846 30096 3851 30152
rect 3734 30092 3740 30094
rect 3804 30092 3851 30096
rect 3785 30091 3851 30092
rect 2576 29952 2896 29953
rect 0 29882 800 29912
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5839 29952 6159 29953
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 29887 6159 29888
rect 9103 29952 9423 29953
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 29887 9423 29888
rect 0 29822 2008 29882
rect 0 29792 800 29822
rect 1948 29746 2008 29822
rect 3877 29746 3943 29749
rect 1948 29744 3943 29746
rect 1948 29688 3882 29744
rect 3938 29688 3943 29744
rect 1948 29686 3943 29688
rect 3877 29683 3943 29686
rect 9489 29474 9555 29477
rect 11200 29474 12000 29504
rect 9489 29472 12000 29474
rect 9489 29416 9494 29472
rect 9550 29416 12000 29472
rect 9489 29414 12000 29416
rect 9489 29411 9555 29414
rect 4207 29408 4527 29409
rect 0 29338 800 29368
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 29343 4527 29344
rect 7471 29408 7791 29409
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 11200 29384 12000 29414
rect 7471 29343 7791 29344
rect 3969 29338 4035 29341
rect 0 29336 4035 29338
rect 0 29280 3974 29336
rect 4030 29280 4035 29336
rect 0 29278 4035 29280
rect 0 29248 800 29278
rect 3969 29275 4035 29278
rect 0 28930 800 28960
rect 0 28870 2514 28930
rect 0 28840 800 28870
rect 2454 28658 2514 28870
rect 2576 28864 2896 28865
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5839 28864 6159 28865
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 28799 6159 28800
rect 9103 28864 9423 28865
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 28799 9423 28800
rect 3141 28796 3207 28797
rect 3141 28794 3188 28796
rect 3096 28792 3188 28794
rect 3096 28736 3146 28792
rect 3096 28734 3188 28736
rect 3141 28732 3188 28734
rect 3252 28732 3258 28796
rect 10133 28794 10199 28797
rect 11200 28794 12000 28824
rect 10133 28792 12000 28794
rect 10133 28736 10138 28792
rect 10194 28736 12000 28792
rect 10133 28734 12000 28736
rect 3141 28731 3207 28732
rect 10133 28731 10199 28734
rect 11200 28704 12000 28734
rect 3233 28658 3299 28661
rect 2454 28656 3299 28658
rect 2454 28600 3238 28656
rect 3294 28600 3299 28656
rect 2454 28598 3299 28600
rect 3233 28595 3299 28598
rect 0 28522 800 28552
rect 2865 28522 2931 28525
rect 0 28520 2931 28522
rect 0 28464 2870 28520
rect 2926 28464 2931 28520
rect 0 28462 2931 28464
rect 0 28432 800 28462
rect 2865 28459 2931 28462
rect 4207 28320 4527 28321
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 28255 4527 28256
rect 7471 28320 7791 28321
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 28255 7791 28256
rect 0 28114 800 28144
rect 1393 28114 1459 28117
rect 0 28112 1459 28114
rect 0 28056 1398 28112
rect 1454 28056 1459 28112
rect 0 28054 1459 28056
rect 0 28024 800 28054
rect 1393 28051 1459 28054
rect 1761 28114 1827 28117
rect 1894 28114 1900 28116
rect 1761 28112 1900 28114
rect 1761 28056 1766 28112
rect 1822 28056 1900 28112
rect 1761 28054 1900 28056
rect 1761 28051 1827 28054
rect 1894 28052 1900 28054
rect 1964 28052 1970 28116
rect 10133 27978 10199 27981
rect 11200 27978 12000 28008
rect 10133 27976 12000 27978
rect 10133 27920 10138 27976
rect 10194 27920 12000 27976
rect 10133 27918 12000 27920
rect 10133 27915 10199 27918
rect 11200 27888 12000 27918
rect 2576 27776 2896 27777
rect 0 27706 800 27736
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5839 27776 6159 27777
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 27711 6159 27712
rect 9103 27776 9423 27777
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 27711 9423 27712
rect 2405 27706 2471 27709
rect 0 27704 2471 27706
rect 0 27648 2410 27704
rect 2466 27648 2471 27704
rect 0 27646 2471 27648
rect 0 27616 800 27646
rect 2405 27643 2471 27646
rect 2037 27570 2103 27573
rect 2998 27570 3004 27572
rect 2037 27568 3004 27570
rect 2037 27512 2042 27568
rect 2098 27512 3004 27568
rect 2037 27510 3004 27512
rect 2037 27507 2103 27510
rect 2998 27508 3004 27510
rect 3068 27508 3074 27572
rect 0 27298 800 27328
rect 2957 27298 3023 27301
rect 0 27296 3023 27298
rect 0 27240 2962 27296
rect 3018 27240 3023 27296
rect 0 27238 3023 27240
rect 0 27208 800 27238
rect 2957 27235 3023 27238
rect 4207 27232 4527 27233
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 27167 4527 27168
rect 7471 27232 7791 27233
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 27167 7791 27168
rect 10133 27162 10199 27165
rect 11200 27162 12000 27192
rect 10133 27160 12000 27162
rect 10133 27104 10138 27160
rect 10194 27104 12000 27160
rect 10133 27102 12000 27104
rect 10133 27099 10199 27102
rect 11200 27072 12000 27102
rect 0 26890 800 26920
rect 3141 26890 3207 26893
rect 0 26888 3207 26890
rect 0 26832 3146 26888
rect 3202 26832 3207 26888
rect 0 26830 3207 26832
rect 0 26800 800 26830
rect 3141 26827 3207 26830
rect 2576 26688 2896 26689
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5839 26688 6159 26689
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 26623 6159 26624
rect 9103 26688 9423 26689
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 26623 9423 26624
rect 10133 26482 10199 26485
rect 11200 26482 12000 26512
rect 10133 26480 12000 26482
rect 10133 26424 10138 26480
rect 10194 26424 12000 26480
rect 10133 26422 12000 26424
rect 10133 26419 10199 26422
rect 11200 26392 12000 26422
rect 0 26346 800 26376
rect 1393 26346 1459 26349
rect 0 26344 1459 26346
rect 0 26288 1398 26344
rect 1454 26288 1459 26344
rect 0 26286 1459 26288
rect 0 26256 800 26286
rect 1393 26283 1459 26286
rect 4207 26144 4527 26145
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 26079 4527 26080
rect 7471 26144 7791 26145
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 26079 7791 26080
rect 0 25938 800 25968
rect 3049 25938 3115 25941
rect 0 25936 3115 25938
rect 0 25880 3054 25936
rect 3110 25880 3115 25936
rect 0 25878 3115 25880
rect 0 25848 800 25878
rect 3049 25875 3115 25878
rect 2865 25802 2931 25805
rect 1488 25800 2931 25802
rect 1488 25744 2870 25800
rect 2926 25744 2931 25800
rect 1488 25742 2931 25744
rect 0 25530 800 25560
rect 1488 25530 1548 25742
rect 2865 25739 2931 25742
rect 10133 25666 10199 25669
rect 11200 25666 12000 25696
rect 10133 25664 12000 25666
rect 10133 25608 10138 25664
rect 10194 25608 12000 25664
rect 10133 25606 12000 25608
rect 10133 25603 10199 25606
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5839 25600 6159 25601
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 25535 6159 25536
rect 9103 25600 9423 25601
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 11200 25576 12000 25606
rect 9103 25535 9423 25536
rect 0 25470 1548 25530
rect 0 25440 800 25470
rect 0 25122 800 25152
rect 1485 25122 1551 25125
rect 0 25120 1551 25122
rect 0 25064 1490 25120
rect 1546 25064 1551 25120
rect 0 25062 1551 25064
rect 0 25032 800 25062
rect 1485 25059 1551 25062
rect 4207 25056 4527 25057
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 24991 4527 24992
rect 7471 25056 7791 25057
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 24991 7791 24992
rect 10133 24850 10199 24853
rect 11200 24850 12000 24880
rect 10133 24848 12000 24850
rect 10133 24792 10138 24848
rect 10194 24792 12000 24848
rect 10133 24790 12000 24792
rect 10133 24787 10199 24790
rect 11200 24760 12000 24790
rect 0 24714 800 24744
rect 2773 24714 2839 24717
rect 0 24712 2839 24714
rect 0 24656 2778 24712
rect 2834 24656 2839 24712
rect 0 24654 2839 24656
rect 0 24624 800 24654
rect 2773 24651 2839 24654
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5839 24512 6159 24513
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 24447 6159 24448
rect 9103 24512 9423 24513
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 24447 9423 24448
rect 0 24306 800 24336
rect 1393 24306 1459 24309
rect 0 24304 1459 24306
rect 0 24248 1398 24304
rect 1454 24248 1459 24304
rect 0 24246 1459 24248
rect 0 24216 800 24246
rect 1393 24243 1459 24246
rect 10133 24170 10199 24173
rect 11200 24170 12000 24200
rect 10133 24168 12000 24170
rect 10133 24112 10138 24168
rect 10194 24112 12000 24168
rect 10133 24110 12000 24112
rect 10133 24107 10199 24110
rect 11200 24080 12000 24110
rect 4207 23968 4527 23969
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 23903 4527 23904
rect 7471 23968 7791 23969
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 23903 7791 23904
rect 0 23762 800 23792
rect 3969 23762 4035 23765
rect 0 23760 4035 23762
rect 0 23704 3974 23760
rect 4030 23704 4035 23760
rect 0 23702 4035 23704
rect 0 23672 800 23702
rect 3969 23699 4035 23702
rect 2576 23424 2896 23425
rect 0 23354 800 23384
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5839 23424 6159 23425
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 23359 6159 23360
rect 9103 23424 9423 23425
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 23359 9423 23360
rect 10041 23354 10107 23357
rect 11200 23354 12000 23384
rect 0 23294 1548 23354
rect 0 23264 800 23294
rect 1488 23218 1548 23294
rect 10041 23352 12000 23354
rect 10041 23296 10046 23352
rect 10102 23296 12000 23352
rect 10041 23294 12000 23296
rect 10041 23291 10107 23294
rect 11200 23264 12000 23294
rect 2957 23218 3023 23221
rect 1488 23216 3023 23218
rect 1488 23160 2962 23216
rect 3018 23160 3023 23216
rect 1488 23158 3023 23160
rect 2957 23155 3023 23158
rect 0 22946 800 22976
rect 1485 22946 1551 22949
rect 0 22944 1551 22946
rect 0 22888 1490 22944
rect 1546 22888 1551 22944
rect 0 22886 1551 22888
rect 0 22856 800 22886
rect 1485 22883 1551 22886
rect 4207 22880 4527 22881
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 22815 4527 22816
rect 7471 22880 7791 22881
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 22815 7791 22816
rect 0 22538 800 22568
rect 3417 22538 3483 22541
rect 0 22536 3483 22538
rect 0 22480 3422 22536
rect 3478 22480 3483 22536
rect 0 22478 3483 22480
rect 0 22448 800 22478
rect 3417 22475 3483 22478
rect 10041 22538 10107 22541
rect 11200 22538 12000 22568
rect 10041 22536 12000 22538
rect 10041 22480 10046 22536
rect 10102 22480 12000 22536
rect 10041 22478 12000 22480
rect 10041 22475 10107 22478
rect 11200 22448 12000 22478
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5839 22336 6159 22337
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 22271 6159 22272
rect 9103 22336 9423 22337
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 22271 9423 22272
rect 0 22130 800 22160
rect 1209 22130 1275 22133
rect 0 22128 1275 22130
rect 0 22072 1214 22128
rect 1270 22072 1275 22128
rect 0 22070 1275 22072
rect 0 22040 800 22070
rect 1209 22067 1275 22070
rect 3182 21932 3188 21996
rect 3252 21994 3258 21996
rect 3601 21994 3667 21997
rect 3252 21992 3667 21994
rect 3252 21936 3606 21992
rect 3662 21936 3667 21992
rect 3252 21934 3667 21936
rect 3252 21932 3258 21934
rect 3601 21931 3667 21934
rect 10041 21858 10107 21861
rect 11200 21858 12000 21888
rect 10041 21856 12000 21858
rect 10041 21800 10046 21856
rect 10102 21800 12000 21856
rect 10041 21798 12000 21800
rect 10041 21795 10107 21798
rect 4207 21792 4527 21793
rect 0 21722 800 21752
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 21727 4527 21728
rect 7471 21792 7791 21793
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 11200 21768 12000 21798
rect 7471 21727 7791 21728
rect 3141 21722 3207 21725
rect 0 21720 3207 21722
rect 0 21664 3146 21720
rect 3202 21664 3207 21720
rect 0 21662 3207 21664
rect 0 21632 800 21662
rect 3141 21659 3207 21662
rect 2576 21248 2896 21249
rect 0 21178 800 21208
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5839 21248 6159 21249
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 21183 6159 21184
rect 9103 21248 9423 21249
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 21183 9423 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 10041 21042 10107 21045
rect 11200 21042 12000 21072
rect 10041 21040 12000 21042
rect 10041 20984 10046 21040
rect 10102 20984 12000 21040
rect 10041 20982 12000 20984
rect 10041 20979 10107 20982
rect 11200 20952 12000 20982
rect 0 20770 800 20800
rect 3969 20770 4035 20773
rect 0 20768 4035 20770
rect 0 20712 3974 20768
rect 4030 20712 4035 20768
rect 0 20710 4035 20712
rect 0 20680 800 20710
rect 3969 20707 4035 20710
rect 4207 20704 4527 20705
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 20639 4527 20640
rect 7471 20704 7791 20705
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 20639 7791 20640
rect 0 20362 800 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 0 20272 800 20302
rect 2773 20299 2839 20302
rect 10041 20362 10107 20365
rect 11200 20362 12000 20392
rect 10041 20360 12000 20362
rect 10041 20304 10046 20360
rect 10102 20304 12000 20360
rect 10041 20302 12000 20304
rect 10041 20299 10107 20302
rect 11200 20272 12000 20302
rect 2576 20160 2896 20161
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5839 20160 6159 20161
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 20095 6159 20096
rect 9103 20160 9423 20161
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 20095 9423 20096
rect 0 19954 800 19984
rect 2957 19954 3023 19957
rect 0 19952 3023 19954
rect 0 19896 2962 19952
rect 3018 19896 3023 19952
rect 0 19894 3023 19896
rect 0 19864 800 19894
rect 2957 19891 3023 19894
rect 4207 19616 4527 19617
rect 0 19546 800 19576
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 19551 4527 19552
rect 7471 19616 7791 19617
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 19551 7791 19552
rect 3141 19546 3207 19549
rect 0 19544 3207 19546
rect 0 19488 3146 19544
rect 3202 19488 3207 19544
rect 0 19486 3207 19488
rect 0 19456 800 19486
rect 3141 19483 3207 19486
rect 10041 19546 10107 19549
rect 11200 19546 12000 19576
rect 10041 19544 12000 19546
rect 10041 19488 10046 19544
rect 10102 19488 12000 19544
rect 10041 19486 12000 19488
rect 10041 19483 10107 19486
rect 11200 19456 12000 19486
rect 2773 19274 2839 19277
rect 1396 19272 2839 19274
rect 1396 19216 2778 19272
rect 2834 19216 2839 19272
rect 1396 19214 2839 19216
rect 0 19138 800 19168
rect 1396 19138 1456 19214
rect 2773 19211 2839 19214
rect 0 19078 1456 19138
rect 0 19048 800 19078
rect 2576 19072 2896 19073
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5839 19072 6159 19073
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 19007 6159 19008
rect 9103 19072 9423 19073
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 19007 9423 19008
rect 10041 18730 10107 18733
rect 11200 18730 12000 18760
rect 10041 18728 12000 18730
rect 10041 18672 10046 18728
rect 10102 18672 12000 18728
rect 10041 18670 12000 18672
rect 10041 18667 10107 18670
rect 11200 18640 12000 18670
rect 0 18594 800 18624
rect 3969 18594 4035 18597
rect 0 18592 4035 18594
rect 0 18536 3974 18592
rect 4030 18536 4035 18592
rect 0 18534 4035 18536
rect 0 18504 800 18534
rect 3969 18531 4035 18534
rect 4207 18528 4527 18529
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 18463 4527 18464
rect 7471 18528 7791 18529
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 18463 7791 18464
rect 0 18186 800 18216
rect 2957 18186 3023 18189
rect 0 18184 3023 18186
rect 0 18128 2962 18184
rect 3018 18128 3023 18184
rect 0 18126 3023 18128
rect 0 18096 800 18126
rect 2957 18123 3023 18126
rect 10041 18050 10107 18053
rect 11200 18050 12000 18080
rect 10041 18048 12000 18050
rect 10041 17992 10046 18048
rect 10102 17992 12000 18048
rect 10041 17990 12000 17992
rect 10041 17987 10107 17990
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5839 17984 6159 17985
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 17919 6159 17920
rect 9103 17984 9423 17985
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 11200 17960 12000 17990
rect 9103 17919 9423 17920
rect 0 17778 800 17808
rect 3417 17778 3483 17781
rect 0 17776 3483 17778
rect 0 17720 3422 17776
rect 3478 17720 3483 17776
rect 0 17718 3483 17720
rect 0 17688 800 17718
rect 3417 17715 3483 17718
rect 4207 17440 4527 17441
rect 0 17370 800 17400
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 17375 4527 17376
rect 7471 17440 7791 17441
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 17375 7791 17376
rect 3969 17370 4035 17373
rect 0 17368 4035 17370
rect 0 17312 3974 17368
rect 4030 17312 4035 17368
rect 0 17310 4035 17312
rect 0 17280 800 17310
rect 3969 17307 4035 17310
rect 10041 17234 10107 17237
rect 11200 17234 12000 17264
rect 10041 17232 12000 17234
rect 10041 17176 10046 17232
rect 10102 17176 12000 17232
rect 10041 17174 12000 17176
rect 10041 17171 10107 17174
rect 11200 17144 12000 17174
rect 2865 17098 2931 17101
rect 1396 17096 2931 17098
rect 1396 17040 2870 17096
rect 2926 17040 2931 17096
rect 1396 17038 2931 17040
rect 0 16962 800 16992
rect 1396 16962 1456 17038
rect 2865 17035 2931 17038
rect 0 16902 1456 16962
rect 0 16872 800 16902
rect 2576 16896 2896 16897
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5839 16896 6159 16897
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 16831 6159 16832
rect 9103 16896 9423 16897
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 16831 9423 16832
rect 0 16554 800 16584
rect 1485 16554 1551 16557
rect 0 16552 1551 16554
rect 0 16496 1490 16552
rect 1546 16496 1551 16552
rect 0 16494 1551 16496
rect 0 16464 800 16494
rect 1485 16491 1551 16494
rect 10041 16418 10107 16421
rect 11200 16418 12000 16448
rect 10041 16416 12000 16418
rect 10041 16360 10046 16416
rect 10102 16360 12000 16416
rect 10041 16358 12000 16360
rect 10041 16355 10107 16358
rect 4207 16352 4527 16353
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 16287 4527 16288
rect 7471 16352 7791 16353
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 11200 16328 12000 16358
rect 7471 16287 7791 16288
rect 0 16010 800 16040
rect 2773 16010 2839 16013
rect 0 16008 2839 16010
rect 0 15952 2778 16008
rect 2834 15952 2839 16008
rect 0 15950 2839 15952
rect 0 15920 800 15950
rect 2773 15947 2839 15950
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5839 15808 6159 15809
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 15743 6159 15744
rect 9103 15808 9423 15809
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 15743 9423 15744
rect 10041 15738 10107 15741
rect 11200 15738 12000 15768
rect 10041 15736 12000 15738
rect 10041 15680 10046 15736
rect 10102 15680 12000 15736
rect 10041 15678 12000 15680
rect 10041 15675 10107 15678
rect 11200 15648 12000 15678
rect 0 15602 800 15632
rect 1393 15602 1459 15605
rect 0 15600 1459 15602
rect 0 15544 1398 15600
rect 1454 15544 1459 15600
rect 0 15542 1459 15544
rect 0 15512 800 15542
rect 1393 15539 1459 15542
rect 4207 15264 4527 15265
rect 0 15194 800 15224
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 15199 4527 15200
rect 7471 15264 7791 15265
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 15199 7791 15200
rect 2865 15194 2931 15197
rect 0 15192 2931 15194
rect 0 15136 2870 15192
rect 2926 15136 2931 15192
rect 0 15134 2931 15136
rect 0 15104 800 15134
rect 2865 15131 2931 15134
rect 10041 14922 10107 14925
rect 11200 14922 12000 14952
rect 10041 14920 12000 14922
rect 10041 14864 10046 14920
rect 10102 14864 12000 14920
rect 10041 14862 12000 14864
rect 10041 14859 10107 14862
rect 11200 14832 12000 14862
rect 0 14786 800 14816
rect 2221 14786 2287 14789
rect 0 14784 2287 14786
rect 0 14728 2226 14784
rect 2282 14728 2287 14784
rect 0 14726 2287 14728
rect 0 14696 800 14726
rect 2221 14723 2287 14726
rect 2576 14720 2896 14721
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5839 14720 6159 14721
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 14655 6159 14656
rect 9103 14720 9423 14721
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 14655 9423 14656
rect 0 14378 800 14408
rect 3969 14378 4035 14381
rect 0 14376 4035 14378
rect 0 14320 3974 14376
rect 4030 14320 4035 14376
rect 0 14318 4035 14320
rect 0 14288 800 14318
rect 3969 14315 4035 14318
rect 4207 14176 4527 14177
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 14111 4527 14112
rect 7471 14176 7791 14177
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 14111 7791 14112
rect 10041 14106 10107 14109
rect 11200 14106 12000 14136
rect 10041 14104 12000 14106
rect 10041 14048 10046 14104
rect 10102 14048 12000 14104
rect 10041 14046 12000 14048
rect 10041 14043 10107 14046
rect 11200 14016 12000 14046
rect 0 13970 800 14000
rect 3141 13970 3207 13973
rect 0 13968 3207 13970
rect 0 13912 3146 13968
rect 3202 13912 3207 13968
rect 0 13910 3207 13912
rect 0 13880 800 13910
rect 3141 13907 3207 13910
rect 2576 13632 2896 13633
rect 0 13562 800 13592
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5839 13632 6159 13633
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 13567 6159 13568
rect 9103 13632 9423 13633
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 13567 9423 13568
rect 1669 13562 1735 13565
rect 0 13560 1735 13562
rect 0 13504 1674 13560
rect 1730 13504 1735 13560
rect 0 13502 1735 13504
rect 0 13472 800 13502
rect 1669 13499 1735 13502
rect 10041 13426 10107 13429
rect 11200 13426 12000 13456
rect 10041 13424 12000 13426
rect 10041 13368 10046 13424
rect 10102 13368 12000 13424
rect 10041 13366 12000 13368
rect 10041 13363 10107 13366
rect 11200 13336 12000 13366
rect 4207 13088 4527 13089
rect 0 13018 800 13048
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 13023 4527 13024
rect 7471 13088 7791 13089
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 13023 7791 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12928 800 12958
rect 2773 12955 2839 12958
rect 0 12610 800 12640
rect 1853 12610 1919 12613
rect 0 12608 1919 12610
rect 0 12552 1858 12608
rect 1914 12552 1919 12608
rect 0 12550 1919 12552
rect 0 12520 800 12550
rect 1853 12547 1919 12550
rect 10041 12610 10107 12613
rect 11200 12610 12000 12640
rect 10041 12608 12000 12610
rect 10041 12552 10046 12608
rect 10102 12552 12000 12608
rect 10041 12550 12000 12552
rect 10041 12547 10107 12550
rect 2576 12544 2896 12545
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5839 12544 6159 12545
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 12479 6159 12480
rect 9103 12544 9423 12545
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 11200 12520 12000 12550
rect 9103 12479 9423 12480
rect 1393 12336 1459 12341
rect 1393 12280 1398 12336
rect 1454 12280 1459 12336
rect 1393 12275 1459 12280
rect 0 12202 800 12232
rect 1396 12202 1456 12275
rect 0 12142 1456 12202
rect 0 12112 800 12142
rect 4207 12000 4527 12001
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 11935 4527 11936
rect 7471 12000 7791 12001
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 11935 7791 11936
rect 0 11794 800 11824
rect 1301 11794 1367 11797
rect 0 11792 1367 11794
rect 0 11736 1306 11792
rect 1362 11736 1367 11792
rect 0 11734 1367 11736
rect 0 11704 800 11734
rect 1301 11731 1367 11734
rect 10041 11794 10107 11797
rect 11200 11794 12000 11824
rect 10041 11792 12000 11794
rect 10041 11736 10046 11792
rect 10102 11736 12000 11792
rect 10041 11734 12000 11736
rect 10041 11731 10107 11734
rect 11200 11704 12000 11734
rect 2576 11456 2896 11457
rect 0 11386 800 11416
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5839 11456 6159 11457
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 11391 6159 11392
rect 9103 11456 9423 11457
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 11391 9423 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 10041 11114 10107 11117
rect 11200 11114 12000 11144
rect 10041 11112 12000 11114
rect 10041 11056 10046 11112
rect 10102 11056 12000 11112
rect 10041 11054 12000 11056
rect 10041 11051 10107 11054
rect 11200 11024 12000 11054
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 4207 10912 4527 10913
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 10847 4527 10848
rect 7471 10912 7791 10913
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 10847 7791 10848
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5839 10368 6159 10369
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 10303 6159 10304
rect 9103 10368 9423 10369
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 10303 9423 10304
rect 10041 10298 10107 10301
rect 11200 10298 12000 10328
rect 10041 10296 12000 10298
rect 10041 10240 10046 10296
rect 10102 10240 12000 10296
rect 10041 10238 12000 10240
rect 10041 10235 10107 10238
rect 11200 10208 12000 10238
rect 0 10026 800 10056
rect 1301 10026 1367 10029
rect 0 10024 1367 10026
rect 0 9968 1306 10024
rect 1362 9968 1367 10024
rect 0 9966 1367 9968
rect 0 9936 800 9966
rect 1301 9963 1367 9966
rect 4207 9824 4527 9825
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 9759 4527 9760
rect 7471 9824 7791 9825
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 9759 7791 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 10041 9482 10107 9485
rect 11200 9482 12000 9512
rect 10041 9480 12000 9482
rect 10041 9424 10046 9480
rect 10102 9424 12000 9480
rect 10041 9422 12000 9424
rect 10041 9419 10107 9422
rect 11200 9392 12000 9422
rect 2576 9280 2896 9281
rect 0 9210 800 9240
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5839 9280 6159 9281
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 9215 6159 9216
rect 9103 9280 9423 9281
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 9215 9423 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 0 8802 800 8832
rect 3049 8802 3115 8805
rect 0 8800 3115 8802
rect 0 8744 3054 8800
rect 3110 8744 3115 8800
rect 0 8742 3115 8744
rect 0 8712 800 8742
rect 3049 8739 3115 8742
rect 10041 8802 10107 8805
rect 11200 8802 12000 8832
rect 10041 8800 12000 8802
rect 10041 8744 10046 8800
rect 10102 8744 12000 8800
rect 10041 8742 12000 8744
rect 10041 8739 10107 8742
rect 4207 8736 4527 8737
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 8671 4527 8672
rect 7471 8736 7791 8737
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 11200 8712 12000 8742
rect 7471 8671 7791 8672
rect 0 8394 800 8424
rect 3509 8394 3575 8397
rect 0 8392 3575 8394
rect 0 8336 3514 8392
rect 3570 8336 3575 8392
rect 0 8334 3575 8336
rect 0 8304 800 8334
rect 3509 8331 3575 8334
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5839 8192 6159 8193
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 8127 6159 8128
rect 9103 8192 9423 8193
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 8127 9423 8128
rect 10041 7986 10107 7989
rect 11200 7986 12000 8016
rect 10041 7984 12000 7986
rect 10041 7928 10046 7984
rect 10102 7928 12000 7984
rect 10041 7926 12000 7928
rect 10041 7923 10107 7926
rect 11200 7896 12000 7926
rect 0 7850 800 7880
rect 3785 7850 3851 7853
rect 0 7848 3851 7850
rect 0 7792 3790 7848
rect 3846 7792 3851 7848
rect 0 7790 3851 7792
rect 0 7760 800 7790
rect 3785 7787 3851 7790
rect 4207 7648 4527 7649
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 7583 4527 7584
rect 7471 7648 7791 7649
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 7583 7791 7584
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 10041 7170 10107 7173
rect 11200 7170 12000 7200
rect 10041 7168 12000 7170
rect 10041 7112 10046 7168
rect 10102 7112 12000 7168
rect 10041 7110 12000 7112
rect 10041 7107 10107 7110
rect 2576 7104 2896 7105
rect 0 7034 800 7064
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5839 7104 6159 7105
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 7039 6159 7040
rect 9103 7104 9423 7105
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 11200 7080 12000 7110
rect 9103 7039 9423 7040
rect 2037 7034 2103 7037
rect 0 7032 2103 7034
rect 0 6976 2042 7032
rect 2098 6976 2103 7032
rect 0 6974 2103 6976
rect 0 6944 800 6974
rect 2037 6971 2103 6974
rect 0 6626 800 6656
rect 1393 6626 1459 6629
rect 0 6624 1459 6626
rect 0 6568 1398 6624
rect 1454 6568 1459 6624
rect 0 6566 1459 6568
rect 0 6536 800 6566
rect 1393 6563 1459 6566
rect 4207 6560 4527 6561
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 6495 4527 6496
rect 7471 6560 7791 6561
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 6495 7791 6496
rect 10041 6490 10107 6493
rect 11200 6490 12000 6520
rect 10041 6488 12000 6490
rect 10041 6432 10046 6488
rect 10102 6432 12000 6488
rect 10041 6430 12000 6432
rect 10041 6427 10107 6430
rect 11200 6400 12000 6430
rect 0 6218 800 6248
rect 3325 6218 3391 6221
rect 0 6216 3391 6218
rect 0 6160 3330 6216
rect 3386 6160 3391 6216
rect 0 6158 3391 6160
rect 0 6128 800 6158
rect 3325 6155 3391 6158
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5839 6016 6159 6017
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 5951 6159 5952
rect 9103 6016 9423 6017
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 5951 9423 5952
rect 0 5810 800 5840
rect 2957 5810 3023 5813
rect 0 5808 3023 5810
rect 0 5752 2962 5808
rect 3018 5752 3023 5808
rect 0 5750 3023 5752
rect 0 5720 800 5750
rect 2957 5747 3023 5750
rect 10041 5674 10107 5677
rect 11200 5674 12000 5704
rect 10041 5672 12000 5674
rect 10041 5616 10046 5672
rect 10102 5616 12000 5672
rect 10041 5614 12000 5616
rect 10041 5611 10107 5614
rect 11200 5584 12000 5614
rect 4207 5472 4527 5473
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 5407 4527 5408
rect 7471 5472 7791 5473
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 5407 7791 5408
rect 0 5266 800 5296
rect 2037 5266 2103 5269
rect 0 5264 2103 5266
rect 0 5208 2042 5264
rect 2098 5208 2103 5264
rect 0 5206 2103 5208
rect 0 5176 800 5206
rect 2037 5203 2103 5206
rect 2576 4928 2896 4929
rect 0 4858 800 4888
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5839 4928 6159 4929
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 4863 6159 4864
rect 9103 4928 9423 4929
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 4863 9423 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 10041 4858 10107 4861
rect 11200 4858 12000 4888
rect 10041 4856 12000 4858
rect 10041 4800 10046 4856
rect 10102 4800 12000 4856
rect 10041 4798 12000 4800
rect 10041 4795 10107 4798
rect 11200 4768 12000 4798
rect 0 4450 800 4480
rect 3969 4450 4035 4453
rect 0 4448 4035 4450
rect 0 4392 3974 4448
rect 4030 4392 4035 4448
rect 0 4390 4035 4392
rect 0 4360 800 4390
rect 3969 4387 4035 4390
rect 4207 4384 4527 4385
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 4319 4527 4320
rect 7471 4384 7791 4385
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 4319 7791 4320
rect 10041 4178 10107 4181
rect 11200 4178 12000 4208
rect 10041 4176 12000 4178
rect 10041 4120 10046 4176
rect 10102 4120 12000 4176
rect 10041 4118 12000 4120
rect 10041 4115 10107 4118
rect 11200 4088 12000 4118
rect 0 4042 800 4072
rect 3969 4042 4035 4045
rect 0 4040 4035 4042
rect 0 3984 3974 4040
rect 4030 3984 4035 4040
rect 0 3982 4035 3984
rect 0 3952 800 3982
rect 3969 3979 4035 3982
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5839 3840 6159 3841
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 3775 6159 3776
rect 9103 3840 9423 3841
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 3775 9423 3776
rect 0 3634 800 3664
rect 1301 3634 1367 3637
rect 0 3632 1367 3634
rect 0 3576 1306 3632
rect 1362 3576 1367 3632
rect 0 3574 1367 3576
rect 0 3544 800 3574
rect 1301 3571 1367 3574
rect 10041 3362 10107 3365
rect 11200 3362 12000 3392
rect 10041 3360 12000 3362
rect 10041 3304 10046 3360
rect 10102 3304 12000 3360
rect 10041 3302 12000 3304
rect 10041 3299 10107 3302
rect 4207 3296 4527 3297
rect 0 3226 800 3256
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 3231 4527 3232
rect 7471 3296 7791 3297
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 11200 3272 12000 3302
rect 7471 3231 7791 3232
rect 1393 3226 1459 3229
rect 0 3224 1459 3226
rect 0 3168 1398 3224
rect 1454 3168 1459 3224
rect 0 3166 1459 3168
rect 0 3136 800 3166
rect 1393 3163 1459 3166
rect 2576 2752 2896 2753
rect 0 2682 800 2712
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5839 2752 6159 2753
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2687 6159 2688
rect 9103 2752 9423 2753
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2687 9423 2688
rect 0 2622 2146 2682
rect 0 2592 800 2622
rect 2086 2546 2146 2622
rect 4061 2546 4127 2549
rect 2086 2544 4127 2546
rect 2086 2488 4066 2544
rect 4122 2488 4127 2544
rect 2086 2486 4127 2488
rect 4061 2483 4127 2486
rect 10041 2546 10107 2549
rect 11200 2546 12000 2576
rect 10041 2544 12000 2546
rect 10041 2488 10046 2544
rect 10102 2488 12000 2544
rect 10041 2486 12000 2488
rect 10041 2483 10107 2486
rect 11200 2456 12000 2486
rect 0 2274 800 2304
rect 3601 2274 3667 2277
rect 0 2272 3667 2274
rect 0 2216 3606 2272
rect 3662 2216 3667 2272
rect 0 2214 3667 2216
rect 0 2184 800 2214
rect 3601 2211 3667 2214
rect 4207 2208 4527 2209
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2143 4527 2144
rect 7471 2208 7791 2209
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2143 7791 2144
rect 0 1866 800 1896
rect 3969 1866 4035 1869
rect 0 1864 4035 1866
rect 0 1808 3974 1864
rect 4030 1808 4035 1864
rect 0 1806 4035 1808
rect 0 1776 800 1806
rect 3969 1803 4035 1806
rect 9489 1866 9555 1869
rect 11200 1866 12000 1896
rect 9489 1864 12000 1866
rect 9489 1808 9494 1864
rect 9550 1808 12000 1864
rect 9489 1806 12000 1808
rect 9489 1803 9555 1806
rect 11200 1776 12000 1806
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 0 1050 800 1080
rect 2865 1050 2931 1053
rect 0 1048 2931 1050
rect 0 992 2870 1048
rect 2926 992 2931 1048
rect 0 990 2931 992
rect 0 960 800 990
rect 2865 987 2931 990
rect 10041 1050 10107 1053
rect 11200 1050 12000 1080
rect 10041 1048 12000 1050
rect 10041 992 10046 1048
rect 10102 992 12000 1048
rect 10041 990 12000 992
rect 10041 987 10107 990
rect 11200 960 12000 990
rect 0 642 800 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 800 582
rect 2773 579 2839 582
rect 9305 370 9371 373
rect 11200 370 12000 400
rect 9305 368 12000 370
rect 9305 312 9310 368
rect 9366 312 12000 368
rect 9305 310 12000 312
rect 9305 307 9371 310
rect 11200 280 12000 310
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5847 77820 5911 77824
rect 5847 77764 5851 77820
rect 5851 77764 5907 77820
rect 5907 77764 5911 77820
rect 5847 77760 5911 77764
rect 5927 77820 5991 77824
rect 5927 77764 5931 77820
rect 5931 77764 5987 77820
rect 5987 77764 5991 77820
rect 5927 77760 5991 77764
rect 6007 77820 6071 77824
rect 6007 77764 6011 77820
rect 6011 77764 6067 77820
rect 6067 77764 6071 77820
rect 6007 77760 6071 77764
rect 6087 77820 6151 77824
rect 6087 77764 6091 77820
rect 6091 77764 6147 77820
rect 6147 77764 6151 77820
rect 6087 77760 6151 77764
rect 9111 77820 9175 77824
rect 9111 77764 9115 77820
rect 9115 77764 9171 77820
rect 9171 77764 9175 77820
rect 9111 77760 9175 77764
rect 9191 77820 9255 77824
rect 9191 77764 9195 77820
rect 9195 77764 9251 77820
rect 9251 77764 9255 77820
rect 9191 77760 9255 77764
rect 9271 77820 9335 77824
rect 9271 77764 9275 77820
rect 9275 77764 9331 77820
rect 9331 77764 9335 77820
rect 9271 77760 9335 77764
rect 9351 77820 9415 77824
rect 9351 77764 9355 77820
rect 9355 77764 9411 77820
rect 9411 77764 9415 77820
rect 9351 77760 9415 77764
rect 4215 77276 4279 77280
rect 4215 77220 4219 77276
rect 4219 77220 4275 77276
rect 4275 77220 4279 77276
rect 4215 77216 4279 77220
rect 4295 77276 4359 77280
rect 4295 77220 4299 77276
rect 4299 77220 4355 77276
rect 4355 77220 4359 77276
rect 4295 77216 4359 77220
rect 4375 77276 4439 77280
rect 4375 77220 4379 77276
rect 4379 77220 4435 77276
rect 4435 77220 4439 77276
rect 4375 77216 4439 77220
rect 4455 77276 4519 77280
rect 4455 77220 4459 77276
rect 4459 77220 4515 77276
rect 4515 77220 4519 77276
rect 4455 77216 4519 77220
rect 7479 77276 7543 77280
rect 7479 77220 7483 77276
rect 7483 77220 7539 77276
rect 7539 77220 7543 77276
rect 7479 77216 7543 77220
rect 7559 77276 7623 77280
rect 7559 77220 7563 77276
rect 7563 77220 7619 77276
rect 7619 77220 7623 77276
rect 7559 77216 7623 77220
rect 7639 77276 7703 77280
rect 7639 77220 7643 77276
rect 7643 77220 7699 77276
rect 7699 77220 7703 77276
rect 7639 77216 7703 77220
rect 7719 77276 7783 77280
rect 7719 77220 7723 77276
rect 7723 77220 7779 77276
rect 7779 77220 7783 77276
rect 7719 77216 7783 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5847 76732 5911 76736
rect 5847 76676 5851 76732
rect 5851 76676 5907 76732
rect 5907 76676 5911 76732
rect 5847 76672 5911 76676
rect 5927 76732 5991 76736
rect 5927 76676 5931 76732
rect 5931 76676 5987 76732
rect 5987 76676 5991 76732
rect 5927 76672 5991 76676
rect 6007 76732 6071 76736
rect 6007 76676 6011 76732
rect 6011 76676 6067 76732
rect 6067 76676 6071 76732
rect 6007 76672 6071 76676
rect 6087 76732 6151 76736
rect 6087 76676 6091 76732
rect 6091 76676 6147 76732
rect 6147 76676 6151 76732
rect 6087 76672 6151 76676
rect 9111 76732 9175 76736
rect 9111 76676 9115 76732
rect 9115 76676 9171 76732
rect 9171 76676 9175 76732
rect 9111 76672 9175 76676
rect 9191 76732 9255 76736
rect 9191 76676 9195 76732
rect 9195 76676 9251 76732
rect 9251 76676 9255 76732
rect 9191 76672 9255 76676
rect 9271 76732 9335 76736
rect 9271 76676 9275 76732
rect 9275 76676 9331 76732
rect 9331 76676 9335 76732
rect 9271 76672 9335 76676
rect 9351 76732 9415 76736
rect 9351 76676 9355 76732
rect 9355 76676 9411 76732
rect 9411 76676 9415 76732
rect 9351 76672 9415 76676
rect 4215 76188 4279 76192
rect 4215 76132 4219 76188
rect 4219 76132 4275 76188
rect 4275 76132 4279 76188
rect 4215 76128 4279 76132
rect 4295 76188 4359 76192
rect 4295 76132 4299 76188
rect 4299 76132 4355 76188
rect 4355 76132 4359 76188
rect 4295 76128 4359 76132
rect 4375 76188 4439 76192
rect 4375 76132 4379 76188
rect 4379 76132 4435 76188
rect 4435 76132 4439 76188
rect 4375 76128 4439 76132
rect 4455 76188 4519 76192
rect 4455 76132 4459 76188
rect 4459 76132 4515 76188
rect 4515 76132 4519 76188
rect 4455 76128 4519 76132
rect 7479 76188 7543 76192
rect 7479 76132 7483 76188
rect 7483 76132 7539 76188
rect 7539 76132 7543 76188
rect 7479 76128 7543 76132
rect 7559 76188 7623 76192
rect 7559 76132 7563 76188
rect 7563 76132 7619 76188
rect 7619 76132 7623 76188
rect 7559 76128 7623 76132
rect 7639 76188 7703 76192
rect 7639 76132 7643 76188
rect 7643 76132 7699 76188
rect 7699 76132 7703 76188
rect 7639 76128 7703 76132
rect 7719 76188 7783 76192
rect 7719 76132 7723 76188
rect 7723 76132 7779 76188
rect 7779 76132 7783 76188
rect 7719 76128 7783 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5847 75644 5911 75648
rect 5847 75588 5851 75644
rect 5851 75588 5907 75644
rect 5907 75588 5911 75644
rect 5847 75584 5911 75588
rect 5927 75644 5991 75648
rect 5927 75588 5931 75644
rect 5931 75588 5987 75644
rect 5987 75588 5991 75644
rect 5927 75584 5991 75588
rect 6007 75644 6071 75648
rect 6007 75588 6011 75644
rect 6011 75588 6067 75644
rect 6067 75588 6071 75644
rect 6007 75584 6071 75588
rect 6087 75644 6151 75648
rect 6087 75588 6091 75644
rect 6091 75588 6147 75644
rect 6147 75588 6151 75644
rect 6087 75584 6151 75588
rect 9111 75644 9175 75648
rect 9111 75588 9115 75644
rect 9115 75588 9171 75644
rect 9171 75588 9175 75644
rect 9111 75584 9175 75588
rect 9191 75644 9255 75648
rect 9191 75588 9195 75644
rect 9195 75588 9251 75644
rect 9251 75588 9255 75644
rect 9191 75584 9255 75588
rect 9271 75644 9335 75648
rect 9271 75588 9275 75644
rect 9275 75588 9331 75644
rect 9331 75588 9335 75644
rect 9271 75584 9335 75588
rect 9351 75644 9415 75648
rect 9351 75588 9355 75644
rect 9355 75588 9411 75644
rect 9411 75588 9415 75644
rect 9351 75584 9415 75588
rect 4215 75100 4279 75104
rect 4215 75044 4219 75100
rect 4219 75044 4275 75100
rect 4275 75044 4279 75100
rect 4215 75040 4279 75044
rect 4295 75100 4359 75104
rect 4295 75044 4299 75100
rect 4299 75044 4355 75100
rect 4355 75044 4359 75100
rect 4295 75040 4359 75044
rect 4375 75100 4439 75104
rect 4375 75044 4379 75100
rect 4379 75044 4435 75100
rect 4435 75044 4439 75100
rect 4375 75040 4439 75044
rect 4455 75100 4519 75104
rect 4455 75044 4459 75100
rect 4459 75044 4515 75100
rect 4515 75044 4519 75100
rect 4455 75040 4519 75044
rect 7479 75100 7543 75104
rect 7479 75044 7483 75100
rect 7483 75044 7539 75100
rect 7539 75044 7543 75100
rect 7479 75040 7543 75044
rect 7559 75100 7623 75104
rect 7559 75044 7563 75100
rect 7563 75044 7619 75100
rect 7619 75044 7623 75100
rect 7559 75040 7623 75044
rect 7639 75100 7703 75104
rect 7639 75044 7643 75100
rect 7643 75044 7699 75100
rect 7699 75044 7703 75100
rect 7639 75040 7703 75044
rect 7719 75100 7783 75104
rect 7719 75044 7723 75100
rect 7723 75044 7779 75100
rect 7779 75044 7783 75100
rect 7719 75040 7783 75044
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5847 74556 5911 74560
rect 5847 74500 5851 74556
rect 5851 74500 5907 74556
rect 5907 74500 5911 74556
rect 5847 74496 5911 74500
rect 5927 74556 5991 74560
rect 5927 74500 5931 74556
rect 5931 74500 5987 74556
rect 5987 74500 5991 74556
rect 5927 74496 5991 74500
rect 6007 74556 6071 74560
rect 6007 74500 6011 74556
rect 6011 74500 6067 74556
rect 6067 74500 6071 74556
rect 6007 74496 6071 74500
rect 6087 74556 6151 74560
rect 6087 74500 6091 74556
rect 6091 74500 6147 74556
rect 6147 74500 6151 74556
rect 6087 74496 6151 74500
rect 9111 74556 9175 74560
rect 9111 74500 9115 74556
rect 9115 74500 9171 74556
rect 9171 74500 9175 74556
rect 9111 74496 9175 74500
rect 9191 74556 9255 74560
rect 9191 74500 9195 74556
rect 9195 74500 9251 74556
rect 9251 74500 9255 74556
rect 9191 74496 9255 74500
rect 9271 74556 9335 74560
rect 9271 74500 9275 74556
rect 9275 74500 9331 74556
rect 9331 74500 9335 74556
rect 9271 74496 9335 74500
rect 9351 74556 9415 74560
rect 9351 74500 9355 74556
rect 9355 74500 9411 74556
rect 9411 74500 9415 74556
rect 9351 74496 9415 74500
rect 4215 74012 4279 74016
rect 4215 73956 4219 74012
rect 4219 73956 4275 74012
rect 4275 73956 4279 74012
rect 4215 73952 4279 73956
rect 4295 74012 4359 74016
rect 4295 73956 4299 74012
rect 4299 73956 4355 74012
rect 4355 73956 4359 74012
rect 4295 73952 4359 73956
rect 4375 74012 4439 74016
rect 4375 73956 4379 74012
rect 4379 73956 4435 74012
rect 4435 73956 4439 74012
rect 4375 73952 4439 73956
rect 4455 74012 4519 74016
rect 4455 73956 4459 74012
rect 4459 73956 4515 74012
rect 4515 73956 4519 74012
rect 4455 73952 4519 73956
rect 7479 74012 7543 74016
rect 7479 73956 7483 74012
rect 7483 73956 7539 74012
rect 7539 73956 7543 74012
rect 7479 73952 7543 73956
rect 7559 74012 7623 74016
rect 7559 73956 7563 74012
rect 7563 73956 7619 74012
rect 7619 73956 7623 74012
rect 7559 73952 7623 73956
rect 7639 74012 7703 74016
rect 7639 73956 7643 74012
rect 7643 73956 7699 74012
rect 7699 73956 7703 74012
rect 7639 73952 7703 73956
rect 7719 74012 7783 74016
rect 7719 73956 7723 74012
rect 7723 73956 7779 74012
rect 7779 73956 7783 74012
rect 7719 73952 7783 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5847 73468 5911 73472
rect 5847 73412 5851 73468
rect 5851 73412 5907 73468
rect 5907 73412 5911 73468
rect 5847 73408 5911 73412
rect 5927 73468 5991 73472
rect 5927 73412 5931 73468
rect 5931 73412 5987 73468
rect 5987 73412 5991 73468
rect 5927 73408 5991 73412
rect 6007 73468 6071 73472
rect 6007 73412 6011 73468
rect 6011 73412 6067 73468
rect 6067 73412 6071 73468
rect 6007 73408 6071 73412
rect 6087 73468 6151 73472
rect 6087 73412 6091 73468
rect 6091 73412 6147 73468
rect 6147 73412 6151 73468
rect 6087 73408 6151 73412
rect 9111 73468 9175 73472
rect 9111 73412 9115 73468
rect 9115 73412 9171 73468
rect 9171 73412 9175 73468
rect 9111 73408 9175 73412
rect 9191 73468 9255 73472
rect 9191 73412 9195 73468
rect 9195 73412 9251 73468
rect 9251 73412 9255 73468
rect 9191 73408 9255 73412
rect 9271 73468 9335 73472
rect 9271 73412 9275 73468
rect 9275 73412 9331 73468
rect 9331 73412 9335 73468
rect 9271 73408 9335 73412
rect 9351 73468 9415 73472
rect 9351 73412 9355 73468
rect 9355 73412 9411 73468
rect 9411 73412 9415 73468
rect 9351 73408 9415 73412
rect 4215 72924 4279 72928
rect 4215 72868 4219 72924
rect 4219 72868 4275 72924
rect 4275 72868 4279 72924
rect 4215 72864 4279 72868
rect 4295 72924 4359 72928
rect 4295 72868 4299 72924
rect 4299 72868 4355 72924
rect 4355 72868 4359 72924
rect 4295 72864 4359 72868
rect 4375 72924 4439 72928
rect 4375 72868 4379 72924
rect 4379 72868 4435 72924
rect 4435 72868 4439 72924
rect 4375 72864 4439 72868
rect 4455 72924 4519 72928
rect 4455 72868 4459 72924
rect 4459 72868 4515 72924
rect 4515 72868 4519 72924
rect 4455 72864 4519 72868
rect 7479 72924 7543 72928
rect 7479 72868 7483 72924
rect 7483 72868 7539 72924
rect 7539 72868 7543 72924
rect 7479 72864 7543 72868
rect 7559 72924 7623 72928
rect 7559 72868 7563 72924
rect 7563 72868 7619 72924
rect 7619 72868 7623 72924
rect 7559 72864 7623 72868
rect 7639 72924 7703 72928
rect 7639 72868 7643 72924
rect 7643 72868 7699 72924
rect 7699 72868 7703 72924
rect 7639 72864 7703 72868
rect 7719 72924 7783 72928
rect 7719 72868 7723 72924
rect 7723 72868 7779 72924
rect 7779 72868 7783 72924
rect 7719 72864 7783 72868
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5847 72380 5911 72384
rect 5847 72324 5851 72380
rect 5851 72324 5907 72380
rect 5907 72324 5911 72380
rect 5847 72320 5911 72324
rect 5927 72380 5991 72384
rect 5927 72324 5931 72380
rect 5931 72324 5987 72380
rect 5987 72324 5991 72380
rect 5927 72320 5991 72324
rect 6007 72380 6071 72384
rect 6007 72324 6011 72380
rect 6011 72324 6067 72380
rect 6067 72324 6071 72380
rect 6007 72320 6071 72324
rect 6087 72380 6151 72384
rect 6087 72324 6091 72380
rect 6091 72324 6147 72380
rect 6147 72324 6151 72380
rect 6087 72320 6151 72324
rect 9111 72380 9175 72384
rect 9111 72324 9115 72380
rect 9115 72324 9171 72380
rect 9171 72324 9175 72380
rect 9111 72320 9175 72324
rect 9191 72380 9255 72384
rect 9191 72324 9195 72380
rect 9195 72324 9251 72380
rect 9251 72324 9255 72380
rect 9191 72320 9255 72324
rect 9271 72380 9335 72384
rect 9271 72324 9275 72380
rect 9275 72324 9331 72380
rect 9331 72324 9335 72380
rect 9271 72320 9335 72324
rect 9351 72380 9415 72384
rect 9351 72324 9355 72380
rect 9355 72324 9411 72380
rect 9411 72324 9415 72380
rect 9351 72320 9415 72324
rect 4215 71836 4279 71840
rect 4215 71780 4219 71836
rect 4219 71780 4275 71836
rect 4275 71780 4279 71836
rect 4215 71776 4279 71780
rect 4295 71836 4359 71840
rect 4295 71780 4299 71836
rect 4299 71780 4355 71836
rect 4355 71780 4359 71836
rect 4295 71776 4359 71780
rect 4375 71836 4439 71840
rect 4375 71780 4379 71836
rect 4379 71780 4435 71836
rect 4435 71780 4439 71836
rect 4375 71776 4439 71780
rect 4455 71836 4519 71840
rect 4455 71780 4459 71836
rect 4459 71780 4515 71836
rect 4515 71780 4519 71836
rect 4455 71776 4519 71780
rect 7479 71836 7543 71840
rect 7479 71780 7483 71836
rect 7483 71780 7539 71836
rect 7539 71780 7543 71836
rect 7479 71776 7543 71780
rect 7559 71836 7623 71840
rect 7559 71780 7563 71836
rect 7563 71780 7619 71836
rect 7619 71780 7623 71836
rect 7559 71776 7623 71780
rect 7639 71836 7703 71840
rect 7639 71780 7643 71836
rect 7643 71780 7699 71836
rect 7699 71780 7703 71836
rect 7639 71776 7703 71780
rect 7719 71836 7783 71840
rect 7719 71780 7723 71836
rect 7723 71780 7779 71836
rect 7779 71780 7783 71836
rect 7719 71776 7783 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5847 71292 5911 71296
rect 5847 71236 5851 71292
rect 5851 71236 5907 71292
rect 5907 71236 5911 71292
rect 5847 71232 5911 71236
rect 5927 71292 5991 71296
rect 5927 71236 5931 71292
rect 5931 71236 5987 71292
rect 5987 71236 5991 71292
rect 5927 71232 5991 71236
rect 6007 71292 6071 71296
rect 6007 71236 6011 71292
rect 6011 71236 6067 71292
rect 6067 71236 6071 71292
rect 6007 71232 6071 71236
rect 6087 71292 6151 71296
rect 6087 71236 6091 71292
rect 6091 71236 6147 71292
rect 6147 71236 6151 71292
rect 6087 71232 6151 71236
rect 9111 71292 9175 71296
rect 9111 71236 9115 71292
rect 9115 71236 9171 71292
rect 9171 71236 9175 71292
rect 9111 71232 9175 71236
rect 9191 71292 9255 71296
rect 9191 71236 9195 71292
rect 9195 71236 9251 71292
rect 9251 71236 9255 71292
rect 9191 71232 9255 71236
rect 9271 71292 9335 71296
rect 9271 71236 9275 71292
rect 9275 71236 9331 71292
rect 9331 71236 9335 71292
rect 9271 71232 9335 71236
rect 9351 71292 9415 71296
rect 9351 71236 9355 71292
rect 9355 71236 9411 71292
rect 9411 71236 9415 71292
rect 9351 71232 9415 71236
rect 4215 70748 4279 70752
rect 4215 70692 4219 70748
rect 4219 70692 4275 70748
rect 4275 70692 4279 70748
rect 4215 70688 4279 70692
rect 4295 70748 4359 70752
rect 4295 70692 4299 70748
rect 4299 70692 4355 70748
rect 4355 70692 4359 70748
rect 4295 70688 4359 70692
rect 4375 70748 4439 70752
rect 4375 70692 4379 70748
rect 4379 70692 4435 70748
rect 4435 70692 4439 70748
rect 4375 70688 4439 70692
rect 4455 70748 4519 70752
rect 4455 70692 4459 70748
rect 4459 70692 4515 70748
rect 4515 70692 4519 70748
rect 4455 70688 4519 70692
rect 7479 70748 7543 70752
rect 7479 70692 7483 70748
rect 7483 70692 7539 70748
rect 7539 70692 7543 70748
rect 7479 70688 7543 70692
rect 7559 70748 7623 70752
rect 7559 70692 7563 70748
rect 7563 70692 7619 70748
rect 7619 70692 7623 70748
rect 7559 70688 7623 70692
rect 7639 70748 7703 70752
rect 7639 70692 7643 70748
rect 7643 70692 7699 70748
rect 7699 70692 7703 70748
rect 7639 70688 7703 70692
rect 7719 70748 7783 70752
rect 7719 70692 7723 70748
rect 7723 70692 7779 70748
rect 7779 70692 7783 70748
rect 7719 70688 7783 70692
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5847 70204 5911 70208
rect 5847 70148 5851 70204
rect 5851 70148 5907 70204
rect 5907 70148 5911 70204
rect 5847 70144 5911 70148
rect 5927 70204 5991 70208
rect 5927 70148 5931 70204
rect 5931 70148 5987 70204
rect 5987 70148 5991 70204
rect 5927 70144 5991 70148
rect 6007 70204 6071 70208
rect 6007 70148 6011 70204
rect 6011 70148 6067 70204
rect 6067 70148 6071 70204
rect 6007 70144 6071 70148
rect 6087 70204 6151 70208
rect 6087 70148 6091 70204
rect 6091 70148 6147 70204
rect 6147 70148 6151 70204
rect 6087 70144 6151 70148
rect 9111 70204 9175 70208
rect 9111 70148 9115 70204
rect 9115 70148 9171 70204
rect 9171 70148 9175 70204
rect 9111 70144 9175 70148
rect 9191 70204 9255 70208
rect 9191 70148 9195 70204
rect 9195 70148 9251 70204
rect 9251 70148 9255 70204
rect 9191 70144 9255 70148
rect 9271 70204 9335 70208
rect 9271 70148 9275 70204
rect 9275 70148 9331 70204
rect 9331 70148 9335 70204
rect 9271 70144 9335 70148
rect 9351 70204 9415 70208
rect 9351 70148 9355 70204
rect 9355 70148 9411 70204
rect 9411 70148 9415 70204
rect 9351 70144 9415 70148
rect 4215 69660 4279 69664
rect 4215 69604 4219 69660
rect 4219 69604 4275 69660
rect 4275 69604 4279 69660
rect 4215 69600 4279 69604
rect 4295 69660 4359 69664
rect 4295 69604 4299 69660
rect 4299 69604 4355 69660
rect 4355 69604 4359 69660
rect 4295 69600 4359 69604
rect 4375 69660 4439 69664
rect 4375 69604 4379 69660
rect 4379 69604 4435 69660
rect 4435 69604 4439 69660
rect 4375 69600 4439 69604
rect 4455 69660 4519 69664
rect 4455 69604 4459 69660
rect 4459 69604 4515 69660
rect 4515 69604 4519 69660
rect 4455 69600 4519 69604
rect 7479 69660 7543 69664
rect 7479 69604 7483 69660
rect 7483 69604 7539 69660
rect 7539 69604 7543 69660
rect 7479 69600 7543 69604
rect 7559 69660 7623 69664
rect 7559 69604 7563 69660
rect 7563 69604 7619 69660
rect 7619 69604 7623 69660
rect 7559 69600 7623 69604
rect 7639 69660 7703 69664
rect 7639 69604 7643 69660
rect 7643 69604 7699 69660
rect 7699 69604 7703 69660
rect 7639 69600 7703 69604
rect 7719 69660 7783 69664
rect 7719 69604 7723 69660
rect 7723 69604 7779 69660
rect 7779 69604 7783 69660
rect 7719 69600 7783 69604
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5847 69116 5911 69120
rect 5847 69060 5851 69116
rect 5851 69060 5907 69116
rect 5907 69060 5911 69116
rect 5847 69056 5911 69060
rect 5927 69116 5991 69120
rect 5927 69060 5931 69116
rect 5931 69060 5987 69116
rect 5987 69060 5991 69116
rect 5927 69056 5991 69060
rect 6007 69116 6071 69120
rect 6007 69060 6011 69116
rect 6011 69060 6067 69116
rect 6067 69060 6071 69116
rect 6007 69056 6071 69060
rect 6087 69116 6151 69120
rect 6087 69060 6091 69116
rect 6091 69060 6147 69116
rect 6147 69060 6151 69116
rect 6087 69056 6151 69060
rect 9111 69116 9175 69120
rect 9111 69060 9115 69116
rect 9115 69060 9171 69116
rect 9171 69060 9175 69116
rect 9111 69056 9175 69060
rect 9191 69116 9255 69120
rect 9191 69060 9195 69116
rect 9195 69060 9251 69116
rect 9251 69060 9255 69116
rect 9191 69056 9255 69060
rect 9271 69116 9335 69120
rect 9271 69060 9275 69116
rect 9275 69060 9331 69116
rect 9331 69060 9335 69116
rect 9271 69056 9335 69060
rect 9351 69116 9415 69120
rect 9351 69060 9355 69116
rect 9355 69060 9411 69116
rect 9411 69060 9415 69116
rect 9351 69056 9415 69060
rect 4215 68572 4279 68576
rect 4215 68516 4219 68572
rect 4219 68516 4275 68572
rect 4275 68516 4279 68572
rect 4215 68512 4279 68516
rect 4295 68572 4359 68576
rect 4295 68516 4299 68572
rect 4299 68516 4355 68572
rect 4355 68516 4359 68572
rect 4295 68512 4359 68516
rect 4375 68572 4439 68576
rect 4375 68516 4379 68572
rect 4379 68516 4435 68572
rect 4435 68516 4439 68572
rect 4375 68512 4439 68516
rect 4455 68572 4519 68576
rect 4455 68516 4459 68572
rect 4459 68516 4515 68572
rect 4515 68516 4519 68572
rect 4455 68512 4519 68516
rect 7479 68572 7543 68576
rect 7479 68516 7483 68572
rect 7483 68516 7539 68572
rect 7539 68516 7543 68572
rect 7479 68512 7543 68516
rect 7559 68572 7623 68576
rect 7559 68516 7563 68572
rect 7563 68516 7619 68572
rect 7619 68516 7623 68572
rect 7559 68512 7623 68516
rect 7639 68572 7703 68576
rect 7639 68516 7643 68572
rect 7643 68516 7699 68572
rect 7699 68516 7703 68572
rect 7639 68512 7703 68516
rect 7719 68572 7783 68576
rect 7719 68516 7723 68572
rect 7723 68516 7779 68572
rect 7779 68516 7783 68572
rect 7719 68512 7783 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5847 68028 5911 68032
rect 5847 67972 5851 68028
rect 5851 67972 5907 68028
rect 5907 67972 5911 68028
rect 5847 67968 5911 67972
rect 5927 68028 5991 68032
rect 5927 67972 5931 68028
rect 5931 67972 5987 68028
rect 5987 67972 5991 68028
rect 5927 67968 5991 67972
rect 6007 68028 6071 68032
rect 6007 67972 6011 68028
rect 6011 67972 6067 68028
rect 6067 67972 6071 68028
rect 6007 67968 6071 67972
rect 6087 68028 6151 68032
rect 6087 67972 6091 68028
rect 6091 67972 6147 68028
rect 6147 67972 6151 68028
rect 6087 67968 6151 67972
rect 9111 68028 9175 68032
rect 9111 67972 9115 68028
rect 9115 67972 9171 68028
rect 9171 67972 9175 68028
rect 9111 67968 9175 67972
rect 9191 68028 9255 68032
rect 9191 67972 9195 68028
rect 9195 67972 9251 68028
rect 9251 67972 9255 68028
rect 9191 67968 9255 67972
rect 9271 68028 9335 68032
rect 9271 67972 9275 68028
rect 9275 67972 9331 68028
rect 9331 67972 9335 68028
rect 9271 67968 9335 67972
rect 9351 68028 9415 68032
rect 9351 67972 9355 68028
rect 9355 67972 9411 68028
rect 9411 67972 9415 68028
rect 9351 67968 9415 67972
rect 4215 67484 4279 67488
rect 4215 67428 4219 67484
rect 4219 67428 4275 67484
rect 4275 67428 4279 67484
rect 4215 67424 4279 67428
rect 4295 67484 4359 67488
rect 4295 67428 4299 67484
rect 4299 67428 4355 67484
rect 4355 67428 4359 67484
rect 4295 67424 4359 67428
rect 4375 67484 4439 67488
rect 4375 67428 4379 67484
rect 4379 67428 4435 67484
rect 4435 67428 4439 67484
rect 4375 67424 4439 67428
rect 4455 67484 4519 67488
rect 4455 67428 4459 67484
rect 4459 67428 4515 67484
rect 4515 67428 4519 67484
rect 4455 67424 4519 67428
rect 7479 67484 7543 67488
rect 7479 67428 7483 67484
rect 7483 67428 7539 67484
rect 7539 67428 7543 67484
rect 7479 67424 7543 67428
rect 7559 67484 7623 67488
rect 7559 67428 7563 67484
rect 7563 67428 7619 67484
rect 7619 67428 7623 67484
rect 7559 67424 7623 67428
rect 7639 67484 7703 67488
rect 7639 67428 7643 67484
rect 7643 67428 7699 67484
rect 7699 67428 7703 67484
rect 7639 67424 7703 67428
rect 7719 67484 7783 67488
rect 7719 67428 7723 67484
rect 7723 67428 7779 67484
rect 7779 67428 7783 67484
rect 7719 67424 7783 67428
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5847 66940 5911 66944
rect 5847 66884 5851 66940
rect 5851 66884 5907 66940
rect 5907 66884 5911 66940
rect 5847 66880 5911 66884
rect 5927 66940 5991 66944
rect 5927 66884 5931 66940
rect 5931 66884 5987 66940
rect 5987 66884 5991 66940
rect 5927 66880 5991 66884
rect 6007 66940 6071 66944
rect 6007 66884 6011 66940
rect 6011 66884 6067 66940
rect 6067 66884 6071 66940
rect 6007 66880 6071 66884
rect 6087 66940 6151 66944
rect 6087 66884 6091 66940
rect 6091 66884 6147 66940
rect 6147 66884 6151 66940
rect 6087 66880 6151 66884
rect 9111 66940 9175 66944
rect 9111 66884 9115 66940
rect 9115 66884 9171 66940
rect 9171 66884 9175 66940
rect 9111 66880 9175 66884
rect 9191 66940 9255 66944
rect 9191 66884 9195 66940
rect 9195 66884 9251 66940
rect 9251 66884 9255 66940
rect 9191 66880 9255 66884
rect 9271 66940 9335 66944
rect 9271 66884 9275 66940
rect 9275 66884 9331 66940
rect 9331 66884 9335 66940
rect 9271 66880 9335 66884
rect 9351 66940 9415 66944
rect 9351 66884 9355 66940
rect 9355 66884 9411 66940
rect 9411 66884 9415 66940
rect 9351 66880 9415 66884
rect 2084 66404 2148 66468
rect 4215 66396 4279 66400
rect 4215 66340 4219 66396
rect 4219 66340 4275 66396
rect 4275 66340 4279 66396
rect 4215 66336 4279 66340
rect 4295 66396 4359 66400
rect 4295 66340 4299 66396
rect 4299 66340 4355 66396
rect 4355 66340 4359 66396
rect 4295 66336 4359 66340
rect 4375 66396 4439 66400
rect 4375 66340 4379 66396
rect 4379 66340 4435 66396
rect 4435 66340 4439 66396
rect 4375 66336 4439 66340
rect 4455 66396 4519 66400
rect 4455 66340 4459 66396
rect 4459 66340 4515 66396
rect 4515 66340 4519 66396
rect 4455 66336 4519 66340
rect 7479 66396 7543 66400
rect 7479 66340 7483 66396
rect 7483 66340 7539 66396
rect 7539 66340 7543 66396
rect 7479 66336 7543 66340
rect 7559 66396 7623 66400
rect 7559 66340 7563 66396
rect 7563 66340 7619 66396
rect 7619 66340 7623 66396
rect 7559 66336 7623 66340
rect 7639 66396 7703 66400
rect 7639 66340 7643 66396
rect 7643 66340 7699 66396
rect 7699 66340 7703 66396
rect 7639 66336 7703 66340
rect 7719 66396 7783 66400
rect 7719 66340 7723 66396
rect 7723 66340 7779 66396
rect 7779 66340 7783 66396
rect 7719 66336 7783 66340
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5847 65852 5911 65856
rect 5847 65796 5851 65852
rect 5851 65796 5907 65852
rect 5907 65796 5911 65852
rect 5847 65792 5911 65796
rect 5927 65852 5991 65856
rect 5927 65796 5931 65852
rect 5931 65796 5987 65852
rect 5987 65796 5991 65852
rect 5927 65792 5991 65796
rect 6007 65852 6071 65856
rect 6007 65796 6011 65852
rect 6011 65796 6067 65852
rect 6067 65796 6071 65852
rect 6007 65792 6071 65796
rect 6087 65852 6151 65856
rect 6087 65796 6091 65852
rect 6091 65796 6147 65852
rect 6147 65796 6151 65852
rect 6087 65792 6151 65796
rect 9111 65852 9175 65856
rect 9111 65796 9115 65852
rect 9115 65796 9171 65852
rect 9171 65796 9175 65852
rect 9111 65792 9175 65796
rect 9191 65852 9255 65856
rect 9191 65796 9195 65852
rect 9195 65796 9251 65852
rect 9251 65796 9255 65852
rect 9191 65792 9255 65796
rect 9271 65852 9335 65856
rect 9271 65796 9275 65852
rect 9275 65796 9331 65852
rect 9331 65796 9335 65852
rect 9271 65792 9335 65796
rect 9351 65852 9415 65856
rect 9351 65796 9355 65852
rect 9355 65796 9411 65852
rect 9411 65796 9415 65852
rect 9351 65792 9415 65796
rect 4215 65308 4279 65312
rect 4215 65252 4219 65308
rect 4219 65252 4275 65308
rect 4275 65252 4279 65308
rect 4215 65248 4279 65252
rect 4295 65308 4359 65312
rect 4295 65252 4299 65308
rect 4299 65252 4355 65308
rect 4355 65252 4359 65308
rect 4295 65248 4359 65252
rect 4375 65308 4439 65312
rect 4375 65252 4379 65308
rect 4379 65252 4435 65308
rect 4435 65252 4439 65308
rect 4375 65248 4439 65252
rect 4455 65308 4519 65312
rect 4455 65252 4459 65308
rect 4459 65252 4515 65308
rect 4515 65252 4519 65308
rect 4455 65248 4519 65252
rect 7479 65308 7543 65312
rect 7479 65252 7483 65308
rect 7483 65252 7539 65308
rect 7539 65252 7543 65308
rect 7479 65248 7543 65252
rect 7559 65308 7623 65312
rect 7559 65252 7563 65308
rect 7563 65252 7619 65308
rect 7619 65252 7623 65308
rect 7559 65248 7623 65252
rect 7639 65308 7703 65312
rect 7639 65252 7643 65308
rect 7643 65252 7699 65308
rect 7699 65252 7703 65308
rect 7639 65248 7703 65252
rect 7719 65308 7783 65312
rect 7719 65252 7723 65308
rect 7723 65252 7779 65308
rect 7779 65252 7783 65308
rect 7719 65248 7783 65252
rect 1900 64908 1964 64972
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5847 64764 5911 64768
rect 5847 64708 5851 64764
rect 5851 64708 5907 64764
rect 5907 64708 5911 64764
rect 5847 64704 5911 64708
rect 5927 64764 5991 64768
rect 5927 64708 5931 64764
rect 5931 64708 5987 64764
rect 5987 64708 5991 64764
rect 5927 64704 5991 64708
rect 6007 64764 6071 64768
rect 6007 64708 6011 64764
rect 6011 64708 6067 64764
rect 6067 64708 6071 64764
rect 6007 64704 6071 64708
rect 6087 64764 6151 64768
rect 6087 64708 6091 64764
rect 6091 64708 6147 64764
rect 6147 64708 6151 64764
rect 6087 64704 6151 64708
rect 9111 64764 9175 64768
rect 9111 64708 9115 64764
rect 9115 64708 9171 64764
rect 9171 64708 9175 64764
rect 9111 64704 9175 64708
rect 9191 64764 9255 64768
rect 9191 64708 9195 64764
rect 9195 64708 9251 64764
rect 9251 64708 9255 64764
rect 9191 64704 9255 64708
rect 9271 64764 9335 64768
rect 9271 64708 9275 64764
rect 9275 64708 9331 64764
rect 9331 64708 9335 64764
rect 9271 64704 9335 64708
rect 9351 64764 9415 64768
rect 9351 64708 9355 64764
rect 9355 64708 9411 64764
rect 9411 64708 9415 64764
rect 9351 64704 9415 64708
rect 4215 64220 4279 64224
rect 4215 64164 4219 64220
rect 4219 64164 4275 64220
rect 4275 64164 4279 64220
rect 4215 64160 4279 64164
rect 4295 64220 4359 64224
rect 4295 64164 4299 64220
rect 4299 64164 4355 64220
rect 4355 64164 4359 64220
rect 4295 64160 4359 64164
rect 4375 64220 4439 64224
rect 4375 64164 4379 64220
rect 4379 64164 4435 64220
rect 4435 64164 4439 64220
rect 4375 64160 4439 64164
rect 4455 64220 4519 64224
rect 4455 64164 4459 64220
rect 4459 64164 4515 64220
rect 4515 64164 4519 64220
rect 4455 64160 4519 64164
rect 7479 64220 7543 64224
rect 7479 64164 7483 64220
rect 7483 64164 7539 64220
rect 7539 64164 7543 64220
rect 7479 64160 7543 64164
rect 7559 64220 7623 64224
rect 7559 64164 7563 64220
rect 7563 64164 7619 64220
rect 7619 64164 7623 64220
rect 7559 64160 7623 64164
rect 7639 64220 7703 64224
rect 7639 64164 7643 64220
rect 7643 64164 7699 64220
rect 7699 64164 7703 64220
rect 7639 64160 7703 64164
rect 7719 64220 7783 64224
rect 7719 64164 7723 64220
rect 7723 64164 7779 64220
rect 7779 64164 7783 64220
rect 7719 64160 7783 64164
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5847 63676 5911 63680
rect 5847 63620 5851 63676
rect 5851 63620 5907 63676
rect 5907 63620 5911 63676
rect 5847 63616 5911 63620
rect 5927 63676 5991 63680
rect 5927 63620 5931 63676
rect 5931 63620 5987 63676
rect 5987 63620 5991 63676
rect 5927 63616 5991 63620
rect 6007 63676 6071 63680
rect 6007 63620 6011 63676
rect 6011 63620 6067 63676
rect 6067 63620 6071 63676
rect 6007 63616 6071 63620
rect 6087 63676 6151 63680
rect 6087 63620 6091 63676
rect 6091 63620 6147 63676
rect 6147 63620 6151 63676
rect 6087 63616 6151 63620
rect 9111 63676 9175 63680
rect 9111 63620 9115 63676
rect 9115 63620 9171 63676
rect 9171 63620 9175 63676
rect 9111 63616 9175 63620
rect 9191 63676 9255 63680
rect 9191 63620 9195 63676
rect 9195 63620 9251 63676
rect 9251 63620 9255 63676
rect 9191 63616 9255 63620
rect 9271 63676 9335 63680
rect 9271 63620 9275 63676
rect 9275 63620 9331 63676
rect 9331 63620 9335 63676
rect 9271 63616 9335 63620
rect 9351 63676 9415 63680
rect 9351 63620 9355 63676
rect 9355 63620 9411 63676
rect 9411 63620 9415 63676
rect 9351 63616 9415 63620
rect 4215 63132 4279 63136
rect 4215 63076 4219 63132
rect 4219 63076 4275 63132
rect 4275 63076 4279 63132
rect 4215 63072 4279 63076
rect 4295 63132 4359 63136
rect 4295 63076 4299 63132
rect 4299 63076 4355 63132
rect 4355 63076 4359 63132
rect 4295 63072 4359 63076
rect 4375 63132 4439 63136
rect 4375 63076 4379 63132
rect 4379 63076 4435 63132
rect 4435 63076 4439 63132
rect 4375 63072 4439 63076
rect 4455 63132 4519 63136
rect 4455 63076 4459 63132
rect 4459 63076 4515 63132
rect 4515 63076 4519 63132
rect 4455 63072 4519 63076
rect 7479 63132 7543 63136
rect 7479 63076 7483 63132
rect 7483 63076 7539 63132
rect 7539 63076 7543 63132
rect 7479 63072 7543 63076
rect 7559 63132 7623 63136
rect 7559 63076 7563 63132
rect 7563 63076 7619 63132
rect 7619 63076 7623 63132
rect 7559 63072 7623 63076
rect 7639 63132 7703 63136
rect 7639 63076 7643 63132
rect 7643 63076 7699 63132
rect 7699 63076 7703 63132
rect 7639 63072 7703 63076
rect 7719 63132 7783 63136
rect 7719 63076 7723 63132
rect 7723 63076 7779 63132
rect 7779 63076 7783 63132
rect 7719 63072 7783 63076
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5847 62588 5911 62592
rect 5847 62532 5851 62588
rect 5851 62532 5907 62588
rect 5907 62532 5911 62588
rect 5847 62528 5911 62532
rect 5927 62588 5991 62592
rect 5927 62532 5931 62588
rect 5931 62532 5987 62588
rect 5987 62532 5991 62588
rect 5927 62528 5991 62532
rect 6007 62588 6071 62592
rect 6007 62532 6011 62588
rect 6011 62532 6067 62588
rect 6067 62532 6071 62588
rect 6007 62528 6071 62532
rect 6087 62588 6151 62592
rect 6087 62532 6091 62588
rect 6091 62532 6147 62588
rect 6147 62532 6151 62588
rect 6087 62528 6151 62532
rect 9111 62588 9175 62592
rect 9111 62532 9115 62588
rect 9115 62532 9171 62588
rect 9171 62532 9175 62588
rect 9111 62528 9175 62532
rect 9191 62588 9255 62592
rect 9191 62532 9195 62588
rect 9195 62532 9251 62588
rect 9251 62532 9255 62588
rect 9191 62528 9255 62532
rect 9271 62588 9335 62592
rect 9271 62532 9275 62588
rect 9275 62532 9331 62588
rect 9331 62532 9335 62588
rect 9271 62528 9335 62532
rect 9351 62588 9415 62592
rect 9351 62532 9355 62588
rect 9355 62532 9411 62588
rect 9411 62532 9415 62588
rect 9351 62528 9415 62532
rect 4215 62044 4279 62048
rect 4215 61988 4219 62044
rect 4219 61988 4275 62044
rect 4275 61988 4279 62044
rect 4215 61984 4279 61988
rect 4295 62044 4359 62048
rect 4295 61988 4299 62044
rect 4299 61988 4355 62044
rect 4355 61988 4359 62044
rect 4295 61984 4359 61988
rect 4375 62044 4439 62048
rect 4375 61988 4379 62044
rect 4379 61988 4435 62044
rect 4435 61988 4439 62044
rect 4375 61984 4439 61988
rect 4455 62044 4519 62048
rect 4455 61988 4459 62044
rect 4459 61988 4515 62044
rect 4515 61988 4519 62044
rect 4455 61984 4519 61988
rect 7479 62044 7543 62048
rect 7479 61988 7483 62044
rect 7483 61988 7539 62044
rect 7539 61988 7543 62044
rect 7479 61984 7543 61988
rect 7559 62044 7623 62048
rect 7559 61988 7563 62044
rect 7563 61988 7619 62044
rect 7619 61988 7623 62044
rect 7559 61984 7623 61988
rect 7639 62044 7703 62048
rect 7639 61988 7643 62044
rect 7643 61988 7699 62044
rect 7699 61988 7703 62044
rect 7639 61984 7703 61988
rect 7719 62044 7783 62048
rect 7719 61988 7723 62044
rect 7723 61988 7779 62044
rect 7779 61988 7783 62044
rect 7719 61984 7783 61988
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5847 61500 5911 61504
rect 5847 61444 5851 61500
rect 5851 61444 5907 61500
rect 5907 61444 5911 61500
rect 5847 61440 5911 61444
rect 5927 61500 5991 61504
rect 5927 61444 5931 61500
rect 5931 61444 5987 61500
rect 5987 61444 5991 61500
rect 5927 61440 5991 61444
rect 6007 61500 6071 61504
rect 6007 61444 6011 61500
rect 6011 61444 6067 61500
rect 6067 61444 6071 61500
rect 6007 61440 6071 61444
rect 6087 61500 6151 61504
rect 6087 61444 6091 61500
rect 6091 61444 6147 61500
rect 6147 61444 6151 61500
rect 6087 61440 6151 61444
rect 9111 61500 9175 61504
rect 9111 61444 9115 61500
rect 9115 61444 9171 61500
rect 9171 61444 9175 61500
rect 9111 61440 9175 61444
rect 9191 61500 9255 61504
rect 9191 61444 9195 61500
rect 9195 61444 9251 61500
rect 9251 61444 9255 61500
rect 9191 61440 9255 61444
rect 9271 61500 9335 61504
rect 9271 61444 9275 61500
rect 9275 61444 9331 61500
rect 9331 61444 9335 61500
rect 9271 61440 9335 61444
rect 9351 61500 9415 61504
rect 9351 61444 9355 61500
rect 9355 61444 9411 61500
rect 9411 61444 9415 61500
rect 9351 61440 9415 61444
rect 4215 60956 4279 60960
rect 4215 60900 4219 60956
rect 4219 60900 4275 60956
rect 4275 60900 4279 60956
rect 4215 60896 4279 60900
rect 4295 60956 4359 60960
rect 4295 60900 4299 60956
rect 4299 60900 4355 60956
rect 4355 60900 4359 60956
rect 4295 60896 4359 60900
rect 4375 60956 4439 60960
rect 4375 60900 4379 60956
rect 4379 60900 4435 60956
rect 4435 60900 4439 60956
rect 4375 60896 4439 60900
rect 4455 60956 4519 60960
rect 4455 60900 4459 60956
rect 4459 60900 4515 60956
rect 4515 60900 4519 60956
rect 4455 60896 4519 60900
rect 7479 60956 7543 60960
rect 7479 60900 7483 60956
rect 7483 60900 7539 60956
rect 7539 60900 7543 60956
rect 7479 60896 7543 60900
rect 7559 60956 7623 60960
rect 7559 60900 7563 60956
rect 7563 60900 7619 60956
rect 7619 60900 7623 60956
rect 7559 60896 7623 60900
rect 7639 60956 7703 60960
rect 7639 60900 7643 60956
rect 7643 60900 7699 60956
rect 7699 60900 7703 60956
rect 7639 60896 7703 60900
rect 7719 60956 7783 60960
rect 7719 60900 7723 60956
rect 7723 60900 7779 60956
rect 7779 60900 7783 60956
rect 7719 60896 7783 60900
rect 2268 60828 2332 60892
rect 2084 60692 2148 60756
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5847 60412 5911 60416
rect 5847 60356 5851 60412
rect 5851 60356 5907 60412
rect 5907 60356 5911 60412
rect 5847 60352 5911 60356
rect 5927 60412 5991 60416
rect 5927 60356 5931 60412
rect 5931 60356 5987 60412
rect 5987 60356 5991 60412
rect 5927 60352 5991 60356
rect 6007 60412 6071 60416
rect 6007 60356 6011 60412
rect 6011 60356 6067 60412
rect 6067 60356 6071 60412
rect 6007 60352 6071 60356
rect 6087 60412 6151 60416
rect 6087 60356 6091 60412
rect 6091 60356 6147 60412
rect 6147 60356 6151 60412
rect 6087 60352 6151 60356
rect 9111 60412 9175 60416
rect 9111 60356 9115 60412
rect 9115 60356 9171 60412
rect 9171 60356 9175 60412
rect 9111 60352 9175 60356
rect 9191 60412 9255 60416
rect 9191 60356 9195 60412
rect 9195 60356 9251 60412
rect 9251 60356 9255 60412
rect 9191 60352 9255 60356
rect 9271 60412 9335 60416
rect 9271 60356 9275 60412
rect 9275 60356 9331 60412
rect 9331 60356 9335 60412
rect 9271 60352 9335 60356
rect 9351 60412 9415 60416
rect 9351 60356 9355 60412
rect 9355 60356 9411 60412
rect 9411 60356 9415 60412
rect 9351 60352 9415 60356
rect 2268 60148 2332 60212
rect 4215 59868 4279 59872
rect 4215 59812 4219 59868
rect 4219 59812 4275 59868
rect 4275 59812 4279 59868
rect 4215 59808 4279 59812
rect 4295 59868 4359 59872
rect 4295 59812 4299 59868
rect 4299 59812 4355 59868
rect 4355 59812 4359 59868
rect 4295 59808 4359 59812
rect 4375 59868 4439 59872
rect 4375 59812 4379 59868
rect 4379 59812 4435 59868
rect 4435 59812 4439 59868
rect 4375 59808 4439 59812
rect 4455 59868 4519 59872
rect 4455 59812 4459 59868
rect 4459 59812 4515 59868
rect 4515 59812 4519 59868
rect 4455 59808 4519 59812
rect 7479 59868 7543 59872
rect 7479 59812 7483 59868
rect 7483 59812 7539 59868
rect 7539 59812 7543 59868
rect 7479 59808 7543 59812
rect 7559 59868 7623 59872
rect 7559 59812 7563 59868
rect 7563 59812 7619 59868
rect 7619 59812 7623 59868
rect 7559 59808 7623 59812
rect 7639 59868 7703 59872
rect 7639 59812 7643 59868
rect 7643 59812 7699 59868
rect 7699 59812 7703 59868
rect 7639 59808 7703 59812
rect 7719 59868 7783 59872
rect 7719 59812 7723 59868
rect 7723 59812 7779 59868
rect 7779 59812 7783 59868
rect 7719 59808 7783 59812
rect 1716 59604 1780 59668
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5847 59324 5911 59328
rect 5847 59268 5851 59324
rect 5851 59268 5907 59324
rect 5907 59268 5911 59324
rect 5847 59264 5911 59268
rect 5927 59324 5991 59328
rect 5927 59268 5931 59324
rect 5931 59268 5987 59324
rect 5987 59268 5991 59324
rect 5927 59264 5991 59268
rect 6007 59324 6071 59328
rect 6007 59268 6011 59324
rect 6011 59268 6067 59324
rect 6067 59268 6071 59324
rect 6007 59264 6071 59268
rect 6087 59324 6151 59328
rect 6087 59268 6091 59324
rect 6091 59268 6147 59324
rect 6147 59268 6151 59324
rect 6087 59264 6151 59268
rect 9111 59324 9175 59328
rect 9111 59268 9115 59324
rect 9115 59268 9171 59324
rect 9171 59268 9175 59324
rect 9111 59264 9175 59268
rect 9191 59324 9255 59328
rect 9191 59268 9195 59324
rect 9195 59268 9251 59324
rect 9251 59268 9255 59324
rect 9191 59264 9255 59268
rect 9271 59324 9335 59328
rect 9271 59268 9275 59324
rect 9275 59268 9331 59324
rect 9331 59268 9335 59324
rect 9271 59264 9335 59268
rect 9351 59324 9415 59328
rect 9351 59268 9355 59324
rect 9355 59268 9411 59324
rect 9411 59268 9415 59324
rect 9351 59264 9415 59268
rect 1900 58788 1964 58852
rect 4215 58780 4279 58784
rect 4215 58724 4219 58780
rect 4219 58724 4275 58780
rect 4275 58724 4279 58780
rect 4215 58720 4279 58724
rect 4295 58780 4359 58784
rect 4295 58724 4299 58780
rect 4299 58724 4355 58780
rect 4355 58724 4359 58780
rect 4295 58720 4359 58724
rect 4375 58780 4439 58784
rect 4375 58724 4379 58780
rect 4379 58724 4435 58780
rect 4435 58724 4439 58780
rect 4375 58720 4439 58724
rect 4455 58780 4519 58784
rect 4455 58724 4459 58780
rect 4459 58724 4515 58780
rect 4515 58724 4519 58780
rect 4455 58720 4519 58724
rect 7479 58780 7543 58784
rect 7479 58724 7483 58780
rect 7483 58724 7539 58780
rect 7539 58724 7543 58780
rect 7479 58720 7543 58724
rect 7559 58780 7623 58784
rect 7559 58724 7563 58780
rect 7563 58724 7619 58780
rect 7619 58724 7623 58780
rect 7559 58720 7623 58724
rect 7639 58780 7703 58784
rect 7639 58724 7643 58780
rect 7643 58724 7699 58780
rect 7699 58724 7703 58780
rect 7639 58720 7703 58724
rect 7719 58780 7783 58784
rect 7719 58724 7723 58780
rect 7723 58724 7779 58780
rect 7779 58724 7783 58780
rect 7719 58720 7783 58724
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5847 58236 5911 58240
rect 5847 58180 5851 58236
rect 5851 58180 5907 58236
rect 5907 58180 5911 58236
rect 5847 58176 5911 58180
rect 5927 58236 5991 58240
rect 5927 58180 5931 58236
rect 5931 58180 5987 58236
rect 5987 58180 5991 58236
rect 5927 58176 5991 58180
rect 6007 58236 6071 58240
rect 6007 58180 6011 58236
rect 6011 58180 6067 58236
rect 6067 58180 6071 58236
rect 6007 58176 6071 58180
rect 6087 58236 6151 58240
rect 6087 58180 6091 58236
rect 6091 58180 6147 58236
rect 6147 58180 6151 58236
rect 6087 58176 6151 58180
rect 9111 58236 9175 58240
rect 9111 58180 9115 58236
rect 9115 58180 9171 58236
rect 9171 58180 9175 58236
rect 9111 58176 9175 58180
rect 9191 58236 9255 58240
rect 9191 58180 9195 58236
rect 9195 58180 9251 58236
rect 9251 58180 9255 58236
rect 9191 58176 9255 58180
rect 9271 58236 9335 58240
rect 9271 58180 9275 58236
rect 9275 58180 9331 58236
rect 9331 58180 9335 58236
rect 9271 58176 9335 58180
rect 9351 58236 9415 58240
rect 9351 58180 9355 58236
rect 9355 58180 9411 58236
rect 9411 58180 9415 58236
rect 9351 58176 9415 58180
rect 3188 57836 3252 57900
rect 4215 57692 4279 57696
rect 4215 57636 4219 57692
rect 4219 57636 4275 57692
rect 4275 57636 4279 57692
rect 4215 57632 4279 57636
rect 4295 57692 4359 57696
rect 4295 57636 4299 57692
rect 4299 57636 4355 57692
rect 4355 57636 4359 57692
rect 4295 57632 4359 57636
rect 4375 57692 4439 57696
rect 4375 57636 4379 57692
rect 4379 57636 4435 57692
rect 4435 57636 4439 57692
rect 4375 57632 4439 57636
rect 4455 57692 4519 57696
rect 4455 57636 4459 57692
rect 4459 57636 4515 57692
rect 4515 57636 4519 57692
rect 4455 57632 4519 57636
rect 7479 57692 7543 57696
rect 7479 57636 7483 57692
rect 7483 57636 7539 57692
rect 7539 57636 7543 57692
rect 7479 57632 7543 57636
rect 7559 57692 7623 57696
rect 7559 57636 7563 57692
rect 7563 57636 7619 57692
rect 7619 57636 7623 57692
rect 7559 57632 7623 57636
rect 7639 57692 7703 57696
rect 7639 57636 7643 57692
rect 7643 57636 7699 57692
rect 7699 57636 7703 57692
rect 7639 57632 7703 57636
rect 7719 57692 7783 57696
rect 7719 57636 7723 57692
rect 7723 57636 7779 57692
rect 7779 57636 7783 57692
rect 7719 57632 7783 57636
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5847 57148 5911 57152
rect 5847 57092 5851 57148
rect 5851 57092 5907 57148
rect 5907 57092 5911 57148
rect 5847 57088 5911 57092
rect 5927 57148 5991 57152
rect 5927 57092 5931 57148
rect 5931 57092 5987 57148
rect 5987 57092 5991 57148
rect 5927 57088 5991 57092
rect 6007 57148 6071 57152
rect 6007 57092 6011 57148
rect 6011 57092 6067 57148
rect 6067 57092 6071 57148
rect 6007 57088 6071 57092
rect 6087 57148 6151 57152
rect 6087 57092 6091 57148
rect 6091 57092 6147 57148
rect 6147 57092 6151 57148
rect 6087 57088 6151 57092
rect 9111 57148 9175 57152
rect 9111 57092 9115 57148
rect 9115 57092 9171 57148
rect 9171 57092 9175 57148
rect 9111 57088 9175 57092
rect 9191 57148 9255 57152
rect 9191 57092 9195 57148
rect 9195 57092 9251 57148
rect 9251 57092 9255 57148
rect 9191 57088 9255 57092
rect 9271 57148 9335 57152
rect 9271 57092 9275 57148
rect 9275 57092 9331 57148
rect 9331 57092 9335 57148
rect 9271 57088 9335 57092
rect 9351 57148 9415 57152
rect 9351 57092 9355 57148
rect 9355 57092 9411 57148
rect 9411 57092 9415 57148
rect 9351 57088 9415 57092
rect 3372 56884 3436 56948
rect 4215 56604 4279 56608
rect 4215 56548 4219 56604
rect 4219 56548 4275 56604
rect 4275 56548 4279 56604
rect 4215 56544 4279 56548
rect 4295 56604 4359 56608
rect 4295 56548 4299 56604
rect 4299 56548 4355 56604
rect 4355 56548 4359 56604
rect 4295 56544 4359 56548
rect 4375 56604 4439 56608
rect 4375 56548 4379 56604
rect 4379 56548 4435 56604
rect 4435 56548 4439 56604
rect 4375 56544 4439 56548
rect 4455 56604 4519 56608
rect 4455 56548 4459 56604
rect 4459 56548 4515 56604
rect 4515 56548 4519 56604
rect 4455 56544 4519 56548
rect 7479 56604 7543 56608
rect 7479 56548 7483 56604
rect 7483 56548 7539 56604
rect 7539 56548 7543 56604
rect 7479 56544 7543 56548
rect 7559 56604 7623 56608
rect 7559 56548 7563 56604
rect 7563 56548 7619 56604
rect 7619 56548 7623 56604
rect 7559 56544 7623 56548
rect 7639 56604 7703 56608
rect 7639 56548 7643 56604
rect 7643 56548 7699 56604
rect 7699 56548 7703 56604
rect 7639 56544 7703 56548
rect 7719 56604 7783 56608
rect 7719 56548 7723 56604
rect 7723 56548 7779 56604
rect 7779 56548 7783 56604
rect 7719 56544 7783 56548
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5847 56060 5911 56064
rect 5847 56004 5851 56060
rect 5851 56004 5907 56060
rect 5907 56004 5911 56060
rect 5847 56000 5911 56004
rect 5927 56060 5991 56064
rect 5927 56004 5931 56060
rect 5931 56004 5987 56060
rect 5987 56004 5991 56060
rect 5927 56000 5991 56004
rect 6007 56060 6071 56064
rect 6007 56004 6011 56060
rect 6011 56004 6067 56060
rect 6067 56004 6071 56060
rect 6007 56000 6071 56004
rect 6087 56060 6151 56064
rect 6087 56004 6091 56060
rect 6091 56004 6147 56060
rect 6147 56004 6151 56060
rect 6087 56000 6151 56004
rect 9111 56060 9175 56064
rect 9111 56004 9115 56060
rect 9115 56004 9171 56060
rect 9171 56004 9175 56060
rect 9111 56000 9175 56004
rect 9191 56060 9255 56064
rect 9191 56004 9195 56060
rect 9195 56004 9251 56060
rect 9251 56004 9255 56060
rect 9191 56000 9255 56004
rect 9271 56060 9335 56064
rect 9271 56004 9275 56060
rect 9275 56004 9331 56060
rect 9331 56004 9335 56060
rect 9271 56000 9335 56004
rect 9351 56060 9415 56064
rect 9351 56004 9355 56060
rect 9355 56004 9411 56060
rect 9411 56004 9415 56060
rect 9351 56000 9415 56004
rect 4215 55516 4279 55520
rect 4215 55460 4219 55516
rect 4219 55460 4275 55516
rect 4275 55460 4279 55516
rect 4215 55456 4279 55460
rect 4295 55516 4359 55520
rect 4295 55460 4299 55516
rect 4299 55460 4355 55516
rect 4355 55460 4359 55516
rect 4295 55456 4359 55460
rect 4375 55516 4439 55520
rect 4375 55460 4379 55516
rect 4379 55460 4435 55516
rect 4435 55460 4439 55516
rect 4375 55456 4439 55460
rect 4455 55516 4519 55520
rect 4455 55460 4459 55516
rect 4459 55460 4515 55516
rect 4515 55460 4519 55516
rect 4455 55456 4519 55460
rect 7479 55516 7543 55520
rect 7479 55460 7483 55516
rect 7483 55460 7539 55516
rect 7539 55460 7543 55516
rect 7479 55456 7543 55460
rect 7559 55516 7623 55520
rect 7559 55460 7563 55516
rect 7563 55460 7619 55516
rect 7619 55460 7623 55516
rect 7559 55456 7623 55460
rect 7639 55516 7703 55520
rect 7639 55460 7643 55516
rect 7643 55460 7699 55516
rect 7699 55460 7703 55516
rect 7639 55456 7703 55460
rect 7719 55516 7783 55520
rect 7719 55460 7723 55516
rect 7723 55460 7779 55516
rect 7779 55460 7783 55516
rect 7719 55456 7783 55460
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 5847 54972 5911 54976
rect 5847 54916 5851 54972
rect 5851 54916 5907 54972
rect 5907 54916 5911 54972
rect 5847 54912 5911 54916
rect 5927 54972 5991 54976
rect 5927 54916 5931 54972
rect 5931 54916 5987 54972
rect 5987 54916 5991 54972
rect 5927 54912 5991 54916
rect 6007 54972 6071 54976
rect 6007 54916 6011 54972
rect 6011 54916 6067 54972
rect 6067 54916 6071 54972
rect 6007 54912 6071 54916
rect 6087 54972 6151 54976
rect 6087 54916 6091 54972
rect 6091 54916 6147 54972
rect 6147 54916 6151 54972
rect 6087 54912 6151 54916
rect 9111 54972 9175 54976
rect 9111 54916 9115 54972
rect 9115 54916 9171 54972
rect 9171 54916 9175 54972
rect 9111 54912 9175 54916
rect 9191 54972 9255 54976
rect 9191 54916 9195 54972
rect 9195 54916 9251 54972
rect 9251 54916 9255 54972
rect 9191 54912 9255 54916
rect 9271 54972 9335 54976
rect 9271 54916 9275 54972
rect 9275 54916 9331 54972
rect 9331 54916 9335 54972
rect 9271 54912 9335 54916
rect 9351 54972 9415 54976
rect 9351 54916 9355 54972
rect 9355 54916 9411 54972
rect 9411 54916 9415 54972
rect 9351 54912 9415 54916
rect 4215 54428 4279 54432
rect 4215 54372 4219 54428
rect 4219 54372 4275 54428
rect 4275 54372 4279 54428
rect 4215 54368 4279 54372
rect 4295 54428 4359 54432
rect 4295 54372 4299 54428
rect 4299 54372 4355 54428
rect 4355 54372 4359 54428
rect 4295 54368 4359 54372
rect 4375 54428 4439 54432
rect 4375 54372 4379 54428
rect 4379 54372 4435 54428
rect 4435 54372 4439 54428
rect 4375 54368 4439 54372
rect 4455 54428 4519 54432
rect 4455 54372 4459 54428
rect 4459 54372 4515 54428
rect 4515 54372 4519 54428
rect 4455 54368 4519 54372
rect 7479 54428 7543 54432
rect 7479 54372 7483 54428
rect 7483 54372 7539 54428
rect 7539 54372 7543 54428
rect 7479 54368 7543 54372
rect 7559 54428 7623 54432
rect 7559 54372 7563 54428
rect 7563 54372 7619 54428
rect 7619 54372 7623 54428
rect 7559 54368 7623 54372
rect 7639 54428 7703 54432
rect 7639 54372 7643 54428
rect 7643 54372 7699 54428
rect 7699 54372 7703 54428
rect 7639 54368 7703 54372
rect 7719 54428 7783 54432
rect 7719 54372 7723 54428
rect 7723 54372 7779 54428
rect 7779 54372 7783 54428
rect 7719 54368 7783 54372
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5847 53884 5911 53888
rect 5847 53828 5851 53884
rect 5851 53828 5907 53884
rect 5907 53828 5911 53884
rect 5847 53824 5911 53828
rect 5927 53884 5991 53888
rect 5927 53828 5931 53884
rect 5931 53828 5987 53884
rect 5987 53828 5991 53884
rect 5927 53824 5991 53828
rect 6007 53884 6071 53888
rect 6007 53828 6011 53884
rect 6011 53828 6067 53884
rect 6067 53828 6071 53884
rect 6007 53824 6071 53828
rect 6087 53884 6151 53888
rect 6087 53828 6091 53884
rect 6091 53828 6147 53884
rect 6147 53828 6151 53884
rect 6087 53824 6151 53828
rect 9111 53884 9175 53888
rect 9111 53828 9115 53884
rect 9115 53828 9171 53884
rect 9171 53828 9175 53884
rect 9111 53824 9175 53828
rect 9191 53884 9255 53888
rect 9191 53828 9195 53884
rect 9195 53828 9251 53884
rect 9251 53828 9255 53884
rect 9191 53824 9255 53828
rect 9271 53884 9335 53888
rect 9271 53828 9275 53884
rect 9275 53828 9331 53884
rect 9331 53828 9335 53884
rect 9271 53824 9335 53828
rect 9351 53884 9415 53888
rect 9351 53828 9355 53884
rect 9355 53828 9411 53884
rect 9411 53828 9415 53884
rect 9351 53824 9415 53828
rect 4215 53340 4279 53344
rect 4215 53284 4219 53340
rect 4219 53284 4275 53340
rect 4275 53284 4279 53340
rect 4215 53280 4279 53284
rect 4295 53340 4359 53344
rect 4295 53284 4299 53340
rect 4299 53284 4355 53340
rect 4355 53284 4359 53340
rect 4295 53280 4359 53284
rect 4375 53340 4439 53344
rect 4375 53284 4379 53340
rect 4379 53284 4435 53340
rect 4435 53284 4439 53340
rect 4375 53280 4439 53284
rect 4455 53340 4519 53344
rect 4455 53284 4459 53340
rect 4459 53284 4515 53340
rect 4515 53284 4519 53340
rect 4455 53280 4519 53284
rect 7479 53340 7543 53344
rect 7479 53284 7483 53340
rect 7483 53284 7539 53340
rect 7539 53284 7543 53340
rect 7479 53280 7543 53284
rect 7559 53340 7623 53344
rect 7559 53284 7563 53340
rect 7563 53284 7619 53340
rect 7619 53284 7623 53340
rect 7559 53280 7623 53284
rect 7639 53340 7703 53344
rect 7639 53284 7643 53340
rect 7643 53284 7699 53340
rect 7699 53284 7703 53340
rect 7639 53280 7703 53284
rect 7719 53340 7783 53344
rect 7719 53284 7723 53340
rect 7723 53284 7779 53340
rect 7779 53284 7783 53340
rect 7719 53280 7783 53284
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5847 52796 5911 52800
rect 5847 52740 5851 52796
rect 5851 52740 5907 52796
rect 5907 52740 5911 52796
rect 5847 52736 5911 52740
rect 5927 52796 5991 52800
rect 5927 52740 5931 52796
rect 5931 52740 5987 52796
rect 5987 52740 5991 52796
rect 5927 52736 5991 52740
rect 6007 52796 6071 52800
rect 6007 52740 6011 52796
rect 6011 52740 6067 52796
rect 6067 52740 6071 52796
rect 6007 52736 6071 52740
rect 6087 52796 6151 52800
rect 6087 52740 6091 52796
rect 6091 52740 6147 52796
rect 6147 52740 6151 52796
rect 6087 52736 6151 52740
rect 9111 52796 9175 52800
rect 9111 52740 9115 52796
rect 9115 52740 9171 52796
rect 9171 52740 9175 52796
rect 9111 52736 9175 52740
rect 9191 52796 9255 52800
rect 9191 52740 9195 52796
rect 9195 52740 9251 52796
rect 9251 52740 9255 52796
rect 9191 52736 9255 52740
rect 9271 52796 9335 52800
rect 9271 52740 9275 52796
rect 9275 52740 9331 52796
rect 9331 52740 9335 52796
rect 9271 52736 9335 52740
rect 9351 52796 9415 52800
rect 9351 52740 9355 52796
rect 9355 52740 9411 52796
rect 9411 52740 9415 52796
rect 9351 52736 9415 52740
rect 4215 52252 4279 52256
rect 4215 52196 4219 52252
rect 4219 52196 4275 52252
rect 4275 52196 4279 52252
rect 4215 52192 4279 52196
rect 4295 52252 4359 52256
rect 4295 52196 4299 52252
rect 4299 52196 4355 52252
rect 4355 52196 4359 52252
rect 4295 52192 4359 52196
rect 4375 52252 4439 52256
rect 4375 52196 4379 52252
rect 4379 52196 4435 52252
rect 4435 52196 4439 52252
rect 4375 52192 4439 52196
rect 4455 52252 4519 52256
rect 4455 52196 4459 52252
rect 4459 52196 4515 52252
rect 4515 52196 4519 52252
rect 4455 52192 4519 52196
rect 7479 52252 7543 52256
rect 7479 52196 7483 52252
rect 7483 52196 7539 52252
rect 7539 52196 7543 52252
rect 7479 52192 7543 52196
rect 7559 52252 7623 52256
rect 7559 52196 7563 52252
rect 7563 52196 7619 52252
rect 7619 52196 7623 52252
rect 7559 52192 7623 52196
rect 7639 52252 7703 52256
rect 7639 52196 7643 52252
rect 7643 52196 7699 52252
rect 7699 52196 7703 52252
rect 7639 52192 7703 52196
rect 7719 52252 7783 52256
rect 7719 52196 7723 52252
rect 7723 52196 7779 52252
rect 7779 52196 7783 52252
rect 7719 52192 7783 52196
rect 1716 51912 1780 51916
rect 1716 51856 1730 51912
rect 1730 51856 1780 51912
rect 1716 51852 1780 51856
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 5847 51708 5911 51712
rect 5847 51652 5851 51708
rect 5851 51652 5907 51708
rect 5907 51652 5911 51708
rect 5847 51648 5911 51652
rect 5927 51708 5991 51712
rect 5927 51652 5931 51708
rect 5931 51652 5987 51708
rect 5987 51652 5991 51708
rect 5927 51648 5991 51652
rect 6007 51708 6071 51712
rect 6007 51652 6011 51708
rect 6011 51652 6067 51708
rect 6067 51652 6071 51708
rect 6007 51648 6071 51652
rect 6087 51708 6151 51712
rect 6087 51652 6091 51708
rect 6091 51652 6147 51708
rect 6147 51652 6151 51708
rect 6087 51648 6151 51652
rect 9111 51708 9175 51712
rect 9111 51652 9115 51708
rect 9115 51652 9171 51708
rect 9171 51652 9175 51708
rect 9111 51648 9175 51652
rect 9191 51708 9255 51712
rect 9191 51652 9195 51708
rect 9195 51652 9251 51708
rect 9251 51652 9255 51708
rect 9191 51648 9255 51652
rect 9271 51708 9335 51712
rect 9271 51652 9275 51708
rect 9275 51652 9331 51708
rect 9331 51652 9335 51708
rect 9271 51648 9335 51652
rect 9351 51708 9415 51712
rect 9351 51652 9355 51708
rect 9355 51652 9411 51708
rect 9411 51652 9415 51708
rect 9351 51648 9415 51652
rect 4215 51164 4279 51168
rect 4215 51108 4219 51164
rect 4219 51108 4275 51164
rect 4275 51108 4279 51164
rect 4215 51104 4279 51108
rect 4295 51164 4359 51168
rect 4295 51108 4299 51164
rect 4299 51108 4355 51164
rect 4355 51108 4359 51164
rect 4295 51104 4359 51108
rect 4375 51164 4439 51168
rect 4375 51108 4379 51164
rect 4379 51108 4435 51164
rect 4435 51108 4439 51164
rect 4375 51104 4439 51108
rect 4455 51164 4519 51168
rect 4455 51108 4459 51164
rect 4459 51108 4515 51164
rect 4515 51108 4519 51164
rect 4455 51104 4519 51108
rect 7479 51164 7543 51168
rect 7479 51108 7483 51164
rect 7483 51108 7539 51164
rect 7539 51108 7543 51164
rect 7479 51104 7543 51108
rect 7559 51164 7623 51168
rect 7559 51108 7563 51164
rect 7563 51108 7619 51164
rect 7619 51108 7623 51164
rect 7559 51104 7623 51108
rect 7639 51164 7703 51168
rect 7639 51108 7643 51164
rect 7643 51108 7699 51164
rect 7699 51108 7703 51164
rect 7639 51104 7703 51108
rect 7719 51164 7783 51168
rect 7719 51108 7723 51164
rect 7723 51108 7779 51164
rect 7779 51108 7783 51164
rect 7719 51104 7783 51108
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5847 50620 5911 50624
rect 5847 50564 5851 50620
rect 5851 50564 5907 50620
rect 5907 50564 5911 50620
rect 5847 50560 5911 50564
rect 5927 50620 5991 50624
rect 5927 50564 5931 50620
rect 5931 50564 5987 50620
rect 5987 50564 5991 50620
rect 5927 50560 5991 50564
rect 6007 50620 6071 50624
rect 6007 50564 6011 50620
rect 6011 50564 6067 50620
rect 6067 50564 6071 50620
rect 6007 50560 6071 50564
rect 6087 50620 6151 50624
rect 6087 50564 6091 50620
rect 6091 50564 6147 50620
rect 6147 50564 6151 50620
rect 6087 50560 6151 50564
rect 9111 50620 9175 50624
rect 9111 50564 9115 50620
rect 9115 50564 9171 50620
rect 9171 50564 9175 50620
rect 9111 50560 9175 50564
rect 9191 50620 9255 50624
rect 9191 50564 9195 50620
rect 9195 50564 9251 50620
rect 9251 50564 9255 50620
rect 9191 50560 9255 50564
rect 9271 50620 9335 50624
rect 9271 50564 9275 50620
rect 9275 50564 9331 50620
rect 9331 50564 9335 50620
rect 9271 50560 9335 50564
rect 9351 50620 9415 50624
rect 9351 50564 9355 50620
rect 9355 50564 9411 50620
rect 9411 50564 9415 50620
rect 9351 50560 9415 50564
rect 3188 50356 3252 50420
rect 4660 50416 4724 50420
rect 4660 50360 4674 50416
rect 4674 50360 4724 50416
rect 4660 50356 4724 50360
rect 4215 50076 4279 50080
rect 4215 50020 4219 50076
rect 4219 50020 4275 50076
rect 4275 50020 4279 50076
rect 4215 50016 4279 50020
rect 4295 50076 4359 50080
rect 4295 50020 4299 50076
rect 4299 50020 4355 50076
rect 4355 50020 4359 50076
rect 4295 50016 4359 50020
rect 4375 50076 4439 50080
rect 4375 50020 4379 50076
rect 4379 50020 4435 50076
rect 4435 50020 4439 50076
rect 4375 50016 4439 50020
rect 4455 50076 4519 50080
rect 4455 50020 4459 50076
rect 4459 50020 4515 50076
rect 4515 50020 4519 50076
rect 4455 50016 4519 50020
rect 7479 50076 7543 50080
rect 7479 50020 7483 50076
rect 7483 50020 7539 50076
rect 7539 50020 7543 50076
rect 7479 50016 7543 50020
rect 7559 50076 7623 50080
rect 7559 50020 7563 50076
rect 7563 50020 7619 50076
rect 7619 50020 7623 50076
rect 7559 50016 7623 50020
rect 7639 50076 7703 50080
rect 7639 50020 7643 50076
rect 7643 50020 7699 50076
rect 7699 50020 7703 50076
rect 7639 50016 7703 50020
rect 7719 50076 7783 50080
rect 7719 50020 7723 50076
rect 7723 50020 7779 50076
rect 7779 50020 7783 50076
rect 7719 50016 7783 50020
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 5847 49532 5911 49536
rect 5847 49476 5851 49532
rect 5851 49476 5907 49532
rect 5907 49476 5911 49532
rect 5847 49472 5911 49476
rect 5927 49532 5991 49536
rect 5927 49476 5931 49532
rect 5931 49476 5987 49532
rect 5987 49476 5991 49532
rect 5927 49472 5991 49476
rect 6007 49532 6071 49536
rect 6007 49476 6011 49532
rect 6011 49476 6067 49532
rect 6067 49476 6071 49532
rect 6007 49472 6071 49476
rect 6087 49532 6151 49536
rect 6087 49476 6091 49532
rect 6091 49476 6147 49532
rect 6147 49476 6151 49532
rect 6087 49472 6151 49476
rect 9111 49532 9175 49536
rect 9111 49476 9115 49532
rect 9115 49476 9171 49532
rect 9171 49476 9175 49532
rect 9111 49472 9175 49476
rect 9191 49532 9255 49536
rect 9191 49476 9195 49532
rect 9195 49476 9251 49532
rect 9251 49476 9255 49532
rect 9191 49472 9255 49476
rect 9271 49532 9335 49536
rect 9271 49476 9275 49532
rect 9275 49476 9331 49532
rect 9331 49476 9335 49532
rect 9271 49472 9335 49476
rect 9351 49532 9415 49536
rect 9351 49476 9355 49532
rect 9355 49476 9411 49532
rect 9411 49476 9415 49532
rect 9351 49472 9415 49476
rect 4215 48988 4279 48992
rect 4215 48932 4219 48988
rect 4219 48932 4275 48988
rect 4275 48932 4279 48988
rect 4215 48928 4279 48932
rect 4295 48988 4359 48992
rect 4295 48932 4299 48988
rect 4299 48932 4355 48988
rect 4355 48932 4359 48988
rect 4295 48928 4359 48932
rect 4375 48988 4439 48992
rect 4375 48932 4379 48988
rect 4379 48932 4435 48988
rect 4435 48932 4439 48988
rect 4375 48928 4439 48932
rect 4455 48988 4519 48992
rect 4455 48932 4459 48988
rect 4459 48932 4515 48988
rect 4515 48932 4519 48988
rect 4455 48928 4519 48932
rect 7479 48988 7543 48992
rect 7479 48932 7483 48988
rect 7483 48932 7539 48988
rect 7539 48932 7543 48988
rect 7479 48928 7543 48932
rect 7559 48988 7623 48992
rect 7559 48932 7563 48988
rect 7563 48932 7619 48988
rect 7619 48932 7623 48988
rect 7559 48928 7623 48932
rect 7639 48988 7703 48992
rect 7639 48932 7643 48988
rect 7643 48932 7699 48988
rect 7699 48932 7703 48988
rect 7639 48928 7703 48932
rect 7719 48988 7783 48992
rect 7719 48932 7723 48988
rect 7723 48932 7779 48988
rect 7779 48932 7783 48988
rect 7719 48928 7783 48932
rect 4660 48724 4724 48788
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 5847 48444 5911 48448
rect 5847 48388 5851 48444
rect 5851 48388 5907 48444
rect 5907 48388 5911 48444
rect 5847 48384 5911 48388
rect 5927 48444 5991 48448
rect 5927 48388 5931 48444
rect 5931 48388 5987 48444
rect 5987 48388 5991 48444
rect 5927 48384 5991 48388
rect 6007 48444 6071 48448
rect 6007 48388 6011 48444
rect 6011 48388 6067 48444
rect 6067 48388 6071 48444
rect 6007 48384 6071 48388
rect 6087 48444 6151 48448
rect 6087 48388 6091 48444
rect 6091 48388 6147 48444
rect 6147 48388 6151 48444
rect 6087 48384 6151 48388
rect 9111 48444 9175 48448
rect 9111 48388 9115 48444
rect 9115 48388 9171 48444
rect 9171 48388 9175 48444
rect 9111 48384 9175 48388
rect 9191 48444 9255 48448
rect 9191 48388 9195 48444
rect 9195 48388 9251 48444
rect 9251 48388 9255 48444
rect 9191 48384 9255 48388
rect 9271 48444 9335 48448
rect 9271 48388 9275 48444
rect 9275 48388 9331 48444
rect 9331 48388 9335 48444
rect 9271 48384 9335 48388
rect 9351 48444 9415 48448
rect 9351 48388 9355 48444
rect 9355 48388 9411 48444
rect 9411 48388 9415 48444
rect 9351 48384 9415 48388
rect 1900 48376 1964 48380
rect 1900 48320 1950 48376
rect 1950 48320 1964 48376
rect 1900 48316 1964 48320
rect 3372 48316 3436 48380
rect 4215 47900 4279 47904
rect 4215 47844 4219 47900
rect 4219 47844 4275 47900
rect 4275 47844 4279 47900
rect 4215 47840 4279 47844
rect 4295 47900 4359 47904
rect 4295 47844 4299 47900
rect 4299 47844 4355 47900
rect 4355 47844 4359 47900
rect 4295 47840 4359 47844
rect 4375 47900 4439 47904
rect 4375 47844 4379 47900
rect 4379 47844 4435 47900
rect 4435 47844 4439 47900
rect 4375 47840 4439 47844
rect 4455 47900 4519 47904
rect 4455 47844 4459 47900
rect 4459 47844 4515 47900
rect 4515 47844 4519 47900
rect 4455 47840 4519 47844
rect 7479 47900 7543 47904
rect 7479 47844 7483 47900
rect 7483 47844 7539 47900
rect 7539 47844 7543 47900
rect 7479 47840 7543 47844
rect 7559 47900 7623 47904
rect 7559 47844 7563 47900
rect 7563 47844 7619 47900
rect 7619 47844 7623 47900
rect 7559 47840 7623 47844
rect 7639 47900 7703 47904
rect 7639 47844 7643 47900
rect 7643 47844 7699 47900
rect 7699 47844 7703 47900
rect 7639 47840 7703 47844
rect 7719 47900 7783 47904
rect 7719 47844 7723 47900
rect 7723 47844 7779 47900
rect 7779 47844 7783 47900
rect 7719 47840 7783 47844
rect 3004 47772 3068 47836
rect 4660 47500 4724 47564
rect 6316 47500 6380 47564
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 5847 47356 5911 47360
rect 5847 47300 5851 47356
rect 5851 47300 5907 47356
rect 5907 47300 5911 47356
rect 5847 47296 5911 47300
rect 5927 47356 5991 47360
rect 5927 47300 5931 47356
rect 5931 47300 5987 47356
rect 5987 47300 5991 47356
rect 5927 47296 5991 47300
rect 6007 47356 6071 47360
rect 6007 47300 6011 47356
rect 6011 47300 6067 47356
rect 6067 47300 6071 47356
rect 6007 47296 6071 47300
rect 6087 47356 6151 47360
rect 6087 47300 6091 47356
rect 6091 47300 6147 47356
rect 6147 47300 6151 47356
rect 6087 47296 6151 47300
rect 9111 47356 9175 47360
rect 9111 47300 9115 47356
rect 9115 47300 9171 47356
rect 9171 47300 9175 47356
rect 9111 47296 9175 47300
rect 9191 47356 9255 47360
rect 9191 47300 9195 47356
rect 9195 47300 9251 47356
rect 9251 47300 9255 47356
rect 9191 47296 9255 47300
rect 9271 47356 9335 47360
rect 9271 47300 9275 47356
rect 9275 47300 9331 47356
rect 9331 47300 9335 47356
rect 9271 47296 9335 47300
rect 9351 47356 9415 47360
rect 9351 47300 9355 47356
rect 9355 47300 9411 47356
rect 9411 47300 9415 47356
rect 9351 47296 9415 47300
rect 2084 47092 2148 47156
rect 4215 46812 4279 46816
rect 4215 46756 4219 46812
rect 4219 46756 4275 46812
rect 4275 46756 4279 46812
rect 4215 46752 4279 46756
rect 4295 46812 4359 46816
rect 4295 46756 4299 46812
rect 4299 46756 4355 46812
rect 4355 46756 4359 46812
rect 4295 46752 4359 46756
rect 4375 46812 4439 46816
rect 4375 46756 4379 46812
rect 4379 46756 4435 46812
rect 4435 46756 4439 46812
rect 4375 46752 4439 46756
rect 4455 46812 4519 46816
rect 4455 46756 4459 46812
rect 4459 46756 4515 46812
rect 4515 46756 4519 46812
rect 4455 46752 4519 46756
rect 7479 46812 7543 46816
rect 7479 46756 7483 46812
rect 7483 46756 7539 46812
rect 7539 46756 7543 46812
rect 7479 46752 7543 46756
rect 7559 46812 7623 46816
rect 7559 46756 7563 46812
rect 7563 46756 7619 46812
rect 7619 46756 7623 46812
rect 7559 46752 7623 46756
rect 7639 46812 7703 46816
rect 7639 46756 7643 46812
rect 7643 46756 7699 46812
rect 7699 46756 7703 46812
rect 7639 46752 7703 46756
rect 7719 46812 7783 46816
rect 7719 46756 7723 46812
rect 7723 46756 7779 46812
rect 7779 46756 7783 46812
rect 7719 46752 7783 46756
rect 3004 46412 3068 46476
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5847 46268 5911 46272
rect 5847 46212 5851 46268
rect 5851 46212 5907 46268
rect 5907 46212 5911 46268
rect 5847 46208 5911 46212
rect 5927 46268 5991 46272
rect 5927 46212 5931 46268
rect 5931 46212 5987 46268
rect 5987 46212 5991 46268
rect 5927 46208 5991 46212
rect 6007 46268 6071 46272
rect 6007 46212 6011 46268
rect 6011 46212 6067 46268
rect 6067 46212 6071 46268
rect 6007 46208 6071 46212
rect 6087 46268 6151 46272
rect 6087 46212 6091 46268
rect 6091 46212 6147 46268
rect 6147 46212 6151 46268
rect 6087 46208 6151 46212
rect 9111 46268 9175 46272
rect 9111 46212 9115 46268
rect 9115 46212 9171 46268
rect 9171 46212 9175 46268
rect 9111 46208 9175 46212
rect 9191 46268 9255 46272
rect 9191 46212 9195 46268
rect 9195 46212 9251 46268
rect 9251 46212 9255 46268
rect 9191 46208 9255 46212
rect 9271 46268 9335 46272
rect 9271 46212 9275 46268
rect 9275 46212 9331 46268
rect 9331 46212 9335 46268
rect 9271 46208 9335 46212
rect 9351 46268 9415 46272
rect 9351 46212 9355 46268
rect 9355 46212 9411 46268
rect 9411 46212 9415 46268
rect 9351 46208 9415 46212
rect 4215 45724 4279 45728
rect 4215 45668 4219 45724
rect 4219 45668 4275 45724
rect 4275 45668 4279 45724
rect 4215 45664 4279 45668
rect 4295 45724 4359 45728
rect 4295 45668 4299 45724
rect 4299 45668 4355 45724
rect 4355 45668 4359 45724
rect 4295 45664 4359 45668
rect 4375 45724 4439 45728
rect 4375 45668 4379 45724
rect 4379 45668 4435 45724
rect 4435 45668 4439 45724
rect 4375 45664 4439 45668
rect 4455 45724 4519 45728
rect 4455 45668 4459 45724
rect 4459 45668 4515 45724
rect 4515 45668 4519 45724
rect 4455 45664 4519 45668
rect 7479 45724 7543 45728
rect 7479 45668 7483 45724
rect 7483 45668 7539 45724
rect 7539 45668 7543 45724
rect 7479 45664 7543 45668
rect 7559 45724 7623 45728
rect 7559 45668 7563 45724
rect 7563 45668 7619 45724
rect 7619 45668 7623 45724
rect 7559 45664 7623 45668
rect 7639 45724 7703 45728
rect 7639 45668 7643 45724
rect 7643 45668 7699 45724
rect 7699 45668 7703 45724
rect 7639 45664 7703 45668
rect 7719 45724 7783 45728
rect 7719 45668 7723 45724
rect 7723 45668 7779 45724
rect 7779 45668 7783 45724
rect 7719 45664 7783 45668
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5847 45180 5911 45184
rect 5847 45124 5851 45180
rect 5851 45124 5907 45180
rect 5907 45124 5911 45180
rect 5847 45120 5911 45124
rect 5927 45180 5991 45184
rect 5927 45124 5931 45180
rect 5931 45124 5987 45180
rect 5987 45124 5991 45180
rect 5927 45120 5991 45124
rect 6007 45180 6071 45184
rect 6007 45124 6011 45180
rect 6011 45124 6067 45180
rect 6067 45124 6071 45180
rect 6007 45120 6071 45124
rect 6087 45180 6151 45184
rect 6087 45124 6091 45180
rect 6091 45124 6147 45180
rect 6147 45124 6151 45180
rect 6087 45120 6151 45124
rect 9111 45180 9175 45184
rect 9111 45124 9115 45180
rect 9115 45124 9171 45180
rect 9171 45124 9175 45180
rect 9111 45120 9175 45124
rect 9191 45180 9255 45184
rect 9191 45124 9195 45180
rect 9195 45124 9251 45180
rect 9251 45124 9255 45180
rect 9191 45120 9255 45124
rect 9271 45180 9335 45184
rect 9271 45124 9275 45180
rect 9275 45124 9331 45180
rect 9331 45124 9335 45180
rect 9271 45120 9335 45124
rect 9351 45180 9415 45184
rect 9351 45124 9355 45180
rect 9355 45124 9411 45180
rect 9411 45124 9415 45180
rect 9351 45120 9415 45124
rect 4215 44636 4279 44640
rect 4215 44580 4219 44636
rect 4219 44580 4275 44636
rect 4275 44580 4279 44636
rect 4215 44576 4279 44580
rect 4295 44636 4359 44640
rect 4295 44580 4299 44636
rect 4299 44580 4355 44636
rect 4355 44580 4359 44636
rect 4295 44576 4359 44580
rect 4375 44636 4439 44640
rect 4375 44580 4379 44636
rect 4379 44580 4435 44636
rect 4435 44580 4439 44636
rect 4375 44576 4439 44580
rect 4455 44636 4519 44640
rect 4455 44580 4459 44636
rect 4459 44580 4515 44636
rect 4515 44580 4519 44636
rect 4455 44576 4519 44580
rect 7479 44636 7543 44640
rect 7479 44580 7483 44636
rect 7483 44580 7539 44636
rect 7539 44580 7543 44636
rect 7479 44576 7543 44580
rect 7559 44636 7623 44640
rect 7559 44580 7563 44636
rect 7563 44580 7619 44636
rect 7619 44580 7623 44636
rect 7559 44576 7623 44580
rect 7639 44636 7703 44640
rect 7639 44580 7643 44636
rect 7643 44580 7699 44636
rect 7699 44580 7703 44636
rect 7639 44576 7703 44580
rect 7719 44636 7783 44640
rect 7719 44580 7723 44636
rect 7723 44580 7779 44636
rect 7779 44580 7783 44636
rect 7719 44576 7783 44580
rect 3004 44372 3068 44436
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5847 44092 5911 44096
rect 5847 44036 5851 44092
rect 5851 44036 5907 44092
rect 5907 44036 5911 44092
rect 5847 44032 5911 44036
rect 5927 44092 5991 44096
rect 5927 44036 5931 44092
rect 5931 44036 5987 44092
rect 5987 44036 5991 44092
rect 5927 44032 5991 44036
rect 6007 44092 6071 44096
rect 6007 44036 6011 44092
rect 6011 44036 6067 44092
rect 6067 44036 6071 44092
rect 6007 44032 6071 44036
rect 6087 44092 6151 44096
rect 6087 44036 6091 44092
rect 6091 44036 6147 44092
rect 6147 44036 6151 44092
rect 6087 44032 6151 44036
rect 9111 44092 9175 44096
rect 9111 44036 9115 44092
rect 9115 44036 9171 44092
rect 9171 44036 9175 44092
rect 9111 44032 9175 44036
rect 9191 44092 9255 44096
rect 9191 44036 9195 44092
rect 9195 44036 9251 44092
rect 9251 44036 9255 44092
rect 9191 44032 9255 44036
rect 9271 44092 9335 44096
rect 9271 44036 9275 44092
rect 9275 44036 9331 44092
rect 9331 44036 9335 44092
rect 9271 44032 9335 44036
rect 9351 44092 9415 44096
rect 9351 44036 9355 44092
rect 9355 44036 9411 44092
rect 9411 44036 9415 44092
rect 9351 44032 9415 44036
rect 6316 43692 6380 43756
rect 4215 43548 4279 43552
rect 4215 43492 4219 43548
rect 4219 43492 4275 43548
rect 4275 43492 4279 43548
rect 4215 43488 4279 43492
rect 4295 43548 4359 43552
rect 4295 43492 4299 43548
rect 4299 43492 4355 43548
rect 4355 43492 4359 43548
rect 4295 43488 4359 43492
rect 4375 43548 4439 43552
rect 4375 43492 4379 43548
rect 4379 43492 4435 43548
rect 4435 43492 4439 43548
rect 4375 43488 4439 43492
rect 4455 43548 4519 43552
rect 4455 43492 4459 43548
rect 4459 43492 4515 43548
rect 4515 43492 4519 43548
rect 4455 43488 4519 43492
rect 7479 43548 7543 43552
rect 7479 43492 7483 43548
rect 7483 43492 7539 43548
rect 7539 43492 7543 43548
rect 7479 43488 7543 43492
rect 7559 43548 7623 43552
rect 7559 43492 7563 43548
rect 7563 43492 7619 43548
rect 7619 43492 7623 43548
rect 7559 43488 7623 43492
rect 7639 43548 7703 43552
rect 7639 43492 7643 43548
rect 7643 43492 7699 43548
rect 7699 43492 7703 43548
rect 7639 43488 7703 43492
rect 7719 43548 7783 43552
rect 7719 43492 7723 43548
rect 7723 43492 7779 43548
rect 7779 43492 7783 43548
rect 7719 43488 7783 43492
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 5847 43004 5911 43008
rect 5847 42948 5851 43004
rect 5851 42948 5907 43004
rect 5907 42948 5911 43004
rect 5847 42944 5911 42948
rect 5927 43004 5991 43008
rect 5927 42948 5931 43004
rect 5931 42948 5987 43004
rect 5987 42948 5991 43004
rect 5927 42944 5991 42948
rect 6007 43004 6071 43008
rect 6007 42948 6011 43004
rect 6011 42948 6067 43004
rect 6067 42948 6071 43004
rect 6007 42944 6071 42948
rect 6087 43004 6151 43008
rect 6087 42948 6091 43004
rect 6091 42948 6147 43004
rect 6147 42948 6151 43004
rect 6087 42944 6151 42948
rect 9111 43004 9175 43008
rect 9111 42948 9115 43004
rect 9115 42948 9171 43004
rect 9171 42948 9175 43004
rect 9111 42944 9175 42948
rect 9191 43004 9255 43008
rect 9191 42948 9195 43004
rect 9195 42948 9251 43004
rect 9251 42948 9255 43004
rect 9191 42944 9255 42948
rect 9271 43004 9335 43008
rect 9271 42948 9275 43004
rect 9275 42948 9331 43004
rect 9331 42948 9335 43004
rect 9271 42944 9335 42948
rect 9351 43004 9415 43008
rect 9351 42948 9355 43004
rect 9355 42948 9411 43004
rect 9411 42948 9415 43004
rect 9351 42944 9415 42948
rect 4660 42468 4724 42532
rect 4215 42460 4279 42464
rect 4215 42404 4219 42460
rect 4219 42404 4275 42460
rect 4275 42404 4279 42460
rect 4215 42400 4279 42404
rect 4295 42460 4359 42464
rect 4295 42404 4299 42460
rect 4299 42404 4355 42460
rect 4355 42404 4359 42460
rect 4295 42400 4359 42404
rect 4375 42460 4439 42464
rect 4375 42404 4379 42460
rect 4379 42404 4435 42460
rect 4435 42404 4439 42460
rect 4375 42400 4439 42404
rect 4455 42460 4519 42464
rect 4455 42404 4459 42460
rect 4459 42404 4515 42460
rect 4515 42404 4519 42460
rect 4455 42400 4519 42404
rect 7479 42460 7543 42464
rect 7479 42404 7483 42460
rect 7483 42404 7539 42460
rect 7539 42404 7543 42460
rect 7479 42400 7543 42404
rect 7559 42460 7623 42464
rect 7559 42404 7563 42460
rect 7563 42404 7619 42460
rect 7619 42404 7623 42460
rect 7559 42400 7623 42404
rect 7639 42460 7703 42464
rect 7639 42404 7643 42460
rect 7643 42404 7699 42460
rect 7699 42404 7703 42460
rect 7639 42400 7703 42404
rect 7719 42460 7783 42464
rect 7719 42404 7723 42460
rect 7723 42404 7779 42460
rect 7779 42404 7783 42460
rect 7719 42400 7783 42404
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5847 41916 5911 41920
rect 5847 41860 5851 41916
rect 5851 41860 5907 41916
rect 5907 41860 5911 41916
rect 5847 41856 5911 41860
rect 5927 41916 5991 41920
rect 5927 41860 5931 41916
rect 5931 41860 5987 41916
rect 5987 41860 5991 41916
rect 5927 41856 5991 41860
rect 6007 41916 6071 41920
rect 6007 41860 6011 41916
rect 6011 41860 6067 41916
rect 6067 41860 6071 41916
rect 6007 41856 6071 41860
rect 6087 41916 6151 41920
rect 6087 41860 6091 41916
rect 6091 41860 6147 41916
rect 6147 41860 6151 41916
rect 6087 41856 6151 41860
rect 9111 41916 9175 41920
rect 9111 41860 9115 41916
rect 9115 41860 9171 41916
rect 9171 41860 9175 41916
rect 9111 41856 9175 41860
rect 9191 41916 9255 41920
rect 9191 41860 9195 41916
rect 9195 41860 9251 41916
rect 9251 41860 9255 41916
rect 9191 41856 9255 41860
rect 9271 41916 9335 41920
rect 9271 41860 9275 41916
rect 9275 41860 9331 41916
rect 9331 41860 9335 41916
rect 9271 41856 9335 41860
rect 9351 41916 9415 41920
rect 9351 41860 9355 41916
rect 9355 41860 9411 41916
rect 9411 41860 9415 41916
rect 9351 41856 9415 41860
rect 3004 41516 3068 41580
rect 4215 41372 4279 41376
rect 4215 41316 4219 41372
rect 4219 41316 4275 41372
rect 4275 41316 4279 41372
rect 4215 41312 4279 41316
rect 4295 41372 4359 41376
rect 4295 41316 4299 41372
rect 4299 41316 4355 41372
rect 4355 41316 4359 41372
rect 4295 41312 4359 41316
rect 4375 41372 4439 41376
rect 4375 41316 4379 41372
rect 4379 41316 4435 41372
rect 4435 41316 4439 41372
rect 4375 41312 4439 41316
rect 4455 41372 4519 41376
rect 4455 41316 4459 41372
rect 4459 41316 4515 41372
rect 4515 41316 4519 41372
rect 4455 41312 4519 41316
rect 7479 41372 7543 41376
rect 7479 41316 7483 41372
rect 7483 41316 7539 41372
rect 7539 41316 7543 41372
rect 7479 41312 7543 41316
rect 7559 41372 7623 41376
rect 7559 41316 7563 41372
rect 7563 41316 7619 41372
rect 7619 41316 7623 41372
rect 7559 41312 7623 41316
rect 7639 41372 7703 41376
rect 7639 41316 7643 41372
rect 7643 41316 7699 41372
rect 7699 41316 7703 41372
rect 7639 41312 7703 41316
rect 7719 41372 7783 41376
rect 7719 41316 7723 41372
rect 7723 41316 7779 41372
rect 7779 41316 7783 41372
rect 7719 41312 7783 41316
rect 2268 41108 2332 41172
rect 3004 41108 3068 41172
rect 2084 40836 2148 40900
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5847 40828 5911 40832
rect 5847 40772 5851 40828
rect 5851 40772 5907 40828
rect 5907 40772 5911 40828
rect 5847 40768 5911 40772
rect 5927 40828 5991 40832
rect 5927 40772 5931 40828
rect 5931 40772 5987 40828
rect 5987 40772 5991 40828
rect 5927 40768 5991 40772
rect 6007 40828 6071 40832
rect 6007 40772 6011 40828
rect 6011 40772 6067 40828
rect 6067 40772 6071 40828
rect 6007 40768 6071 40772
rect 6087 40828 6151 40832
rect 6087 40772 6091 40828
rect 6091 40772 6147 40828
rect 6147 40772 6151 40828
rect 6087 40768 6151 40772
rect 9111 40828 9175 40832
rect 9111 40772 9115 40828
rect 9115 40772 9171 40828
rect 9171 40772 9175 40828
rect 9111 40768 9175 40772
rect 9191 40828 9255 40832
rect 9191 40772 9195 40828
rect 9195 40772 9251 40828
rect 9251 40772 9255 40828
rect 9191 40768 9255 40772
rect 9271 40828 9335 40832
rect 9271 40772 9275 40828
rect 9275 40772 9331 40828
rect 9331 40772 9335 40828
rect 9271 40768 9335 40772
rect 9351 40828 9415 40832
rect 9351 40772 9355 40828
rect 9355 40772 9411 40828
rect 9411 40772 9415 40828
rect 9351 40768 9415 40772
rect 4215 40284 4279 40288
rect 4215 40228 4219 40284
rect 4219 40228 4275 40284
rect 4275 40228 4279 40284
rect 4215 40224 4279 40228
rect 4295 40284 4359 40288
rect 4295 40228 4299 40284
rect 4299 40228 4355 40284
rect 4355 40228 4359 40284
rect 4295 40224 4359 40228
rect 4375 40284 4439 40288
rect 4375 40228 4379 40284
rect 4379 40228 4435 40284
rect 4435 40228 4439 40284
rect 4375 40224 4439 40228
rect 4455 40284 4519 40288
rect 4455 40228 4459 40284
rect 4459 40228 4515 40284
rect 4515 40228 4519 40284
rect 4455 40224 4519 40228
rect 7479 40284 7543 40288
rect 7479 40228 7483 40284
rect 7483 40228 7539 40284
rect 7539 40228 7543 40284
rect 7479 40224 7543 40228
rect 7559 40284 7623 40288
rect 7559 40228 7563 40284
rect 7563 40228 7619 40284
rect 7619 40228 7623 40284
rect 7559 40224 7623 40228
rect 7639 40284 7703 40288
rect 7639 40228 7643 40284
rect 7643 40228 7699 40284
rect 7699 40228 7703 40284
rect 7639 40224 7703 40228
rect 7719 40284 7783 40288
rect 7719 40228 7723 40284
rect 7723 40228 7779 40284
rect 7779 40228 7783 40284
rect 7719 40224 7783 40228
rect 1900 40020 1964 40084
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5847 39740 5911 39744
rect 5847 39684 5851 39740
rect 5851 39684 5907 39740
rect 5907 39684 5911 39740
rect 5847 39680 5911 39684
rect 5927 39740 5991 39744
rect 5927 39684 5931 39740
rect 5931 39684 5987 39740
rect 5987 39684 5991 39740
rect 5927 39680 5991 39684
rect 6007 39740 6071 39744
rect 6007 39684 6011 39740
rect 6011 39684 6067 39740
rect 6067 39684 6071 39740
rect 6007 39680 6071 39684
rect 6087 39740 6151 39744
rect 6087 39684 6091 39740
rect 6091 39684 6147 39740
rect 6147 39684 6151 39740
rect 6087 39680 6151 39684
rect 9111 39740 9175 39744
rect 9111 39684 9115 39740
rect 9115 39684 9171 39740
rect 9171 39684 9175 39740
rect 9111 39680 9175 39684
rect 9191 39740 9255 39744
rect 9191 39684 9195 39740
rect 9195 39684 9251 39740
rect 9251 39684 9255 39740
rect 9191 39680 9255 39684
rect 9271 39740 9335 39744
rect 9271 39684 9275 39740
rect 9275 39684 9331 39740
rect 9331 39684 9335 39740
rect 9271 39680 9335 39684
rect 9351 39740 9415 39744
rect 9351 39684 9355 39740
rect 9355 39684 9411 39740
rect 9411 39684 9415 39740
rect 9351 39680 9415 39684
rect 4215 39196 4279 39200
rect 4215 39140 4219 39196
rect 4219 39140 4275 39196
rect 4275 39140 4279 39196
rect 4215 39136 4279 39140
rect 4295 39196 4359 39200
rect 4295 39140 4299 39196
rect 4299 39140 4355 39196
rect 4355 39140 4359 39196
rect 4295 39136 4359 39140
rect 4375 39196 4439 39200
rect 4375 39140 4379 39196
rect 4379 39140 4435 39196
rect 4435 39140 4439 39196
rect 4375 39136 4439 39140
rect 4455 39196 4519 39200
rect 4455 39140 4459 39196
rect 4459 39140 4515 39196
rect 4515 39140 4519 39196
rect 4455 39136 4519 39140
rect 7479 39196 7543 39200
rect 7479 39140 7483 39196
rect 7483 39140 7539 39196
rect 7539 39140 7543 39196
rect 7479 39136 7543 39140
rect 7559 39196 7623 39200
rect 7559 39140 7563 39196
rect 7563 39140 7619 39196
rect 7619 39140 7623 39196
rect 7559 39136 7623 39140
rect 7639 39196 7703 39200
rect 7639 39140 7643 39196
rect 7643 39140 7699 39196
rect 7699 39140 7703 39196
rect 7639 39136 7703 39140
rect 7719 39196 7783 39200
rect 7719 39140 7723 39196
rect 7723 39140 7779 39196
rect 7779 39140 7783 39196
rect 7719 39136 7783 39140
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5847 38652 5911 38656
rect 5847 38596 5851 38652
rect 5851 38596 5907 38652
rect 5907 38596 5911 38652
rect 5847 38592 5911 38596
rect 5927 38652 5991 38656
rect 5927 38596 5931 38652
rect 5931 38596 5987 38652
rect 5987 38596 5991 38652
rect 5927 38592 5991 38596
rect 6007 38652 6071 38656
rect 6007 38596 6011 38652
rect 6011 38596 6067 38652
rect 6067 38596 6071 38652
rect 6007 38592 6071 38596
rect 6087 38652 6151 38656
rect 6087 38596 6091 38652
rect 6091 38596 6147 38652
rect 6147 38596 6151 38652
rect 6087 38592 6151 38596
rect 9111 38652 9175 38656
rect 9111 38596 9115 38652
rect 9115 38596 9171 38652
rect 9171 38596 9175 38652
rect 9111 38592 9175 38596
rect 9191 38652 9255 38656
rect 9191 38596 9195 38652
rect 9195 38596 9251 38652
rect 9251 38596 9255 38652
rect 9191 38592 9255 38596
rect 9271 38652 9335 38656
rect 9271 38596 9275 38652
rect 9275 38596 9331 38652
rect 9331 38596 9335 38652
rect 9271 38592 9335 38596
rect 9351 38652 9415 38656
rect 9351 38596 9355 38652
rect 9355 38596 9411 38652
rect 9411 38596 9415 38652
rect 9351 38592 9415 38596
rect 3740 38252 3804 38316
rect 4215 38108 4279 38112
rect 4215 38052 4219 38108
rect 4219 38052 4275 38108
rect 4275 38052 4279 38108
rect 4215 38048 4279 38052
rect 4295 38108 4359 38112
rect 4295 38052 4299 38108
rect 4299 38052 4355 38108
rect 4355 38052 4359 38108
rect 4295 38048 4359 38052
rect 4375 38108 4439 38112
rect 4375 38052 4379 38108
rect 4379 38052 4435 38108
rect 4435 38052 4439 38108
rect 4375 38048 4439 38052
rect 4455 38108 4519 38112
rect 4455 38052 4459 38108
rect 4459 38052 4515 38108
rect 4515 38052 4519 38108
rect 4455 38048 4519 38052
rect 7479 38108 7543 38112
rect 7479 38052 7483 38108
rect 7483 38052 7539 38108
rect 7539 38052 7543 38108
rect 7479 38048 7543 38052
rect 7559 38108 7623 38112
rect 7559 38052 7563 38108
rect 7563 38052 7619 38108
rect 7619 38052 7623 38108
rect 7559 38048 7623 38052
rect 7639 38108 7703 38112
rect 7639 38052 7643 38108
rect 7643 38052 7699 38108
rect 7699 38052 7703 38108
rect 7639 38048 7703 38052
rect 7719 38108 7783 38112
rect 7719 38052 7723 38108
rect 7723 38052 7779 38108
rect 7779 38052 7783 38108
rect 7719 38048 7783 38052
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5847 37564 5911 37568
rect 5847 37508 5851 37564
rect 5851 37508 5907 37564
rect 5907 37508 5911 37564
rect 5847 37504 5911 37508
rect 5927 37564 5991 37568
rect 5927 37508 5931 37564
rect 5931 37508 5987 37564
rect 5987 37508 5991 37564
rect 5927 37504 5991 37508
rect 6007 37564 6071 37568
rect 6007 37508 6011 37564
rect 6011 37508 6067 37564
rect 6067 37508 6071 37564
rect 6007 37504 6071 37508
rect 6087 37564 6151 37568
rect 6087 37508 6091 37564
rect 6091 37508 6147 37564
rect 6147 37508 6151 37564
rect 6087 37504 6151 37508
rect 9111 37564 9175 37568
rect 9111 37508 9115 37564
rect 9115 37508 9171 37564
rect 9171 37508 9175 37564
rect 9111 37504 9175 37508
rect 9191 37564 9255 37568
rect 9191 37508 9195 37564
rect 9195 37508 9251 37564
rect 9251 37508 9255 37564
rect 9191 37504 9255 37508
rect 9271 37564 9335 37568
rect 9271 37508 9275 37564
rect 9275 37508 9331 37564
rect 9331 37508 9335 37564
rect 9271 37504 9335 37508
rect 9351 37564 9415 37568
rect 9351 37508 9355 37564
rect 9355 37508 9411 37564
rect 9411 37508 9415 37564
rect 9351 37504 9415 37508
rect 3372 37300 3436 37364
rect 4215 37020 4279 37024
rect 4215 36964 4219 37020
rect 4219 36964 4275 37020
rect 4275 36964 4279 37020
rect 4215 36960 4279 36964
rect 4295 37020 4359 37024
rect 4295 36964 4299 37020
rect 4299 36964 4355 37020
rect 4355 36964 4359 37020
rect 4295 36960 4359 36964
rect 4375 37020 4439 37024
rect 4375 36964 4379 37020
rect 4379 36964 4435 37020
rect 4435 36964 4439 37020
rect 4375 36960 4439 36964
rect 4455 37020 4519 37024
rect 4455 36964 4459 37020
rect 4459 36964 4515 37020
rect 4515 36964 4519 37020
rect 4455 36960 4519 36964
rect 7479 37020 7543 37024
rect 7479 36964 7483 37020
rect 7483 36964 7539 37020
rect 7539 36964 7543 37020
rect 7479 36960 7543 36964
rect 7559 37020 7623 37024
rect 7559 36964 7563 37020
rect 7563 36964 7619 37020
rect 7619 36964 7623 37020
rect 7559 36960 7623 36964
rect 7639 37020 7703 37024
rect 7639 36964 7643 37020
rect 7643 36964 7699 37020
rect 7699 36964 7703 37020
rect 7639 36960 7703 36964
rect 7719 37020 7783 37024
rect 7719 36964 7723 37020
rect 7723 36964 7779 37020
rect 7779 36964 7783 37020
rect 7719 36960 7783 36964
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5847 36476 5911 36480
rect 5847 36420 5851 36476
rect 5851 36420 5907 36476
rect 5907 36420 5911 36476
rect 5847 36416 5911 36420
rect 5927 36476 5991 36480
rect 5927 36420 5931 36476
rect 5931 36420 5987 36476
rect 5987 36420 5991 36476
rect 5927 36416 5991 36420
rect 6007 36476 6071 36480
rect 6007 36420 6011 36476
rect 6011 36420 6067 36476
rect 6067 36420 6071 36476
rect 6007 36416 6071 36420
rect 6087 36476 6151 36480
rect 6087 36420 6091 36476
rect 6091 36420 6147 36476
rect 6147 36420 6151 36476
rect 6087 36416 6151 36420
rect 9111 36476 9175 36480
rect 9111 36420 9115 36476
rect 9115 36420 9171 36476
rect 9171 36420 9175 36476
rect 9111 36416 9175 36420
rect 9191 36476 9255 36480
rect 9191 36420 9195 36476
rect 9195 36420 9251 36476
rect 9251 36420 9255 36476
rect 9191 36416 9255 36420
rect 9271 36476 9335 36480
rect 9271 36420 9275 36476
rect 9275 36420 9331 36476
rect 9331 36420 9335 36476
rect 9271 36416 9335 36420
rect 9351 36476 9415 36480
rect 9351 36420 9355 36476
rect 9355 36420 9411 36476
rect 9411 36420 9415 36476
rect 9351 36416 9415 36420
rect 4215 35932 4279 35936
rect 4215 35876 4219 35932
rect 4219 35876 4275 35932
rect 4275 35876 4279 35932
rect 4215 35872 4279 35876
rect 4295 35932 4359 35936
rect 4295 35876 4299 35932
rect 4299 35876 4355 35932
rect 4355 35876 4359 35932
rect 4295 35872 4359 35876
rect 4375 35932 4439 35936
rect 4375 35876 4379 35932
rect 4379 35876 4435 35932
rect 4435 35876 4439 35932
rect 4375 35872 4439 35876
rect 4455 35932 4519 35936
rect 4455 35876 4459 35932
rect 4459 35876 4515 35932
rect 4515 35876 4519 35932
rect 4455 35872 4519 35876
rect 7479 35932 7543 35936
rect 7479 35876 7483 35932
rect 7483 35876 7539 35932
rect 7539 35876 7543 35932
rect 7479 35872 7543 35876
rect 7559 35932 7623 35936
rect 7559 35876 7563 35932
rect 7563 35876 7619 35932
rect 7619 35876 7623 35932
rect 7559 35872 7623 35876
rect 7639 35932 7703 35936
rect 7639 35876 7643 35932
rect 7643 35876 7699 35932
rect 7699 35876 7703 35932
rect 7639 35872 7703 35876
rect 7719 35932 7783 35936
rect 7719 35876 7723 35932
rect 7723 35876 7779 35932
rect 7779 35876 7783 35932
rect 7719 35872 7783 35876
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5847 35388 5911 35392
rect 5847 35332 5851 35388
rect 5851 35332 5907 35388
rect 5907 35332 5911 35388
rect 5847 35328 5911 35332
rect 5927 35388 5991 35392
rect 5927 35332 5931 35388
rect 5931 35332 5987 35388
rect 5987 35332 5991 35388
rect 5927 35328 5991 35332
rect 6007 35388 6071 35392
rect 6007 35332 6011 35388
rect 6011 35332 6067 35388
rect 6067 35332 6071 35388
rect 6007 35328 6071 35332
rect 6087 35388 6151 35392
rect 6087 35332 6091 35388
rect 6091 35332 6147 35388
rect 6147 35332 6151 35388
rect 6087 35328 6151 35332
rect 9111 35388 9175 35392
rect 9111 35332 9115 35388
rect 9115 35332 9171 35388
rect 9171 35332 9175 35388
rect 9111 35328 9175 35332
rect 9191 35388 9255 35392
rect 9191 35332 9195 35388
rect 9195 35332 9251 35388
rect 9251 35332 9255 35388
rect 9191 35328 9255 35332
rect 9271 35388 9335 35392
rect 9271 35332 9275 35388
rect 9275 35332 9331 35388
rect 9331 35332 9335 35388
rect 9271 35328 9335 35332
rect 9351 35388 9415 35392
rect 9351 35332 9355 35388
rect 9355 35332 9411 35388
rect 9411 35332 9415 35388
rect 9351 35328 9415 35332
rect 4215 34844 4279 34848
rect 4215 34788 4219 34844
rect 4219 34788 4275 34844
rect 4275 34788 4279 34844
rect 4215 34784 4279 34788
rect 4295 34844 4359 34848
rect 4295 34788 4299 34844
rect 4299 34788 4355 34844
rect 4355 34788 4359 34844
rect 4295 34784 4359 34788
rect 4375 34844 4439 34848
rect 4375 34788 4379 34844
rect 4379 34788 4435 34844
rect 4435 34788 4439 34844
rect 4375 34784 4439 34788
rect 4455 34844 4519 34848
rect 4455 34788 4459 34844
rect 4459 34788 4515 34844
rect 4515 34788 4519 34844
rect 4455 34784 4519 34788
rect 7479 34844 7543 34848
rect 7479 34788 7483 34844
rect 7483 34788 7539 34844
rect 7539 34788 7543 34844
rect 7479 34784 7543 34788
rect 7559 34844 7623 34848
rect 7559 34788 7563 34844
rect 7563 34788 7619 34844
rect 7619 34788 7623 34844
rect 7559 34784 7623 34788
rect 7639 34844 7703 34848
rect 7639 34788 7643 34844
rect 7643 34788 7699 34844
rect 7699 34788 7703 34844
rect 7639 34784 7703 34788
rect 7719 34844 7783 34848
rect 7719 34788 7723 34844
rect 7723 34788 7779 34844
rect 7779 34788 7783 34844
rect 7719 34784 7783 34788
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5847 34300 5911 34304
rect 5847 34244 5851 34300
rect 5851 34244 5907 34300
rect 5907 34244 5911 34300
rect 5847 34240 5911 34244
rect 5927 34300 5991 34304
rect 5927 34244 5931 34300
rect 5931 34244 5987 34300
rect 5987 34244 5991 34300
rect 5927 34240 5991 34244
rect 6007 34300 6071 34304
rect 6007 34244 6011 34300
rect 6011 34244 6067 34300
rect 6067 34244 6071 34300
rect 6007 34240 6071 34244
rect 6087 34300 6151 34304
rect 6087 34244 6091 34300
rect 6091 34244 6147 34300
rect 6147 34244 6151 34300
rect 6087 34240 6151 34244
rect 9111 34300 9175 34304
rect 9111 34244 9115 34300
rect 9115 34244 9171 34300
rect 9171 34244 9175 34300
rect 9111 34240 9175 34244
rect 9191 34300 9255 34304
rect 9191 34244 9195 34300
rect 9195 34244 9251 34300
rect 9251 34244 9255 34300
rect 9191 34240 9255 34244
rect 9271 34300 9335 34304
rect 9271 34244 9275 34300
rect 9275 34244 9331 34300
rect 9331 34244 9335 34300
rect 9271 34240 9335 34244
rect 9351 34300 9415 34304
rect 9351 34244 9355 34300
rect 9355 34244 9411 34300
rect 9411 34244 9415 34300
rect 9351 34240 9415 34244
rect 4215 33756 4279 33760
rect 4215 33700 4219 33756
rect 4219 33700 4275 33756
rect 4275 33700 4279 33756
rect 4215 33696 4279 33700
rect 4295 33756 4359 33760
rect 4295 33700 4299 33756
rect 4299 33700 4355 33756
rect 4355 33700 4359 33756
rect 4295 33696 4359 33700
rect 4375 33756 4439 33760
rect 4375 33700 4379 33756
rect 4379 33700 4435 33756
rect 4435 33700 4439 33756
rect 4375 33696 4439 33700
rect 4455 33756 4519 33760
rect 4455 33700 4459 33756
rect 4459 33700 4515 33756
rect 4515 33700 4519 33756
rect 4455 33696 4519 33700
rect 7479 33756 7543 33760
rect 7479 33700 7483 33756
rect 7483 33700 7539 33756
rect 7539 33700 7543 33756
rect 7479 33696 7543 33700
rect 7559 33756 7623 33760
rect 7559 33700 7563 33756
rect 7563 33700 7619 33756
rect 7619 33700 7623 33756
rect 7559 33696 7623 33700
rect 7639 33756 7703 33760
rect 7639 33700 7643 33756
rect 7643 33700 7699 33756
rect 7699 33700 7703 33756
rect 7639 33696 7703 33700
rect 7719 33756 7783 33760
rect 7719 33700 7723 33756
rect 7723 33700 7779 33756
rect 7779 33700 7783 33756
rect 7719 33696 7783 33700
rect 3372 33492 3436 33556
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5847 33212 5911 33216
rect 5847 33156 5851 33212
rect 5851 33156 5907 33212
rect 5907 33156 5911 33212
rect 5847 33152 5911 33156
rect 5927 33212 5991 33216
rect 5927 33156 5931 33212
rect 5931 33156 5987 33212
rect 5987 33156 5991 33212
rect 5927 33152 5991 33156
rect 6007 33212 6071 33216
rect 6007 33156 6011 33212
rect 6011 33156 6067 33212
rect 6067 33156 6071 33212
rect 6007 33152 6071 33156
rect 6087 33212 6151 33216
rect 6087 33156 6091 33212
rect 6091 33156 6147 33212
rect 6147 33156 6151 33212
rect 6087 33152 6151 33156
rect 9111 33212 9175 33216
rect 9111 33156 9115 33212
rect 9115 33156 9171 33212
rect 9171 33156 9175 33212
rect 9111 33152 9175 33156
rect 9191 33212 9255 33216
rect 9191 33156 9195 33212
rect 9195 33156 9251 33212
rect 9251 33156 9255 33212
rect 9191 33152 9255 33156
rect 9271 33212 9335 33216
rect 9271 33156 9275 33212
rect 9275 33156 9331 33212
rect 9331 33156 9335 33212
rect 9271 33152 9335 33156
rect 9351 33212 9415 33216
rect 9351 33156 9355 33212
rect 9355 33156 9411 33212
rect 9411 33156 9415 33212
rect 9351 33152 9415 33156
rect 4215 32668 4279 32672
rect 4215 32612 4219 32668
rect 4219 32612 4275 32668
rect 4275 32612 4279 32668
rect 4215 32608 4279 32612
rect 4295 32668 4359 32672
rect 4295 32612 4299 32668
rect 4299 32612 4355 32668
rect 4355 32612 4359 32668
rect 4295 32608 4359 32612
rect 4375 32668 4439 32672
rect 4375 32612 4379 32668
rect 4379 32612 4435 32668
rect 4435 32612 4439 32668
rect 4375 32608 4439 32612
rect 4455 32668 4519 32672
rect 4455 32612 4459 32668
rect 4459 32612 4515 32668
rect 4515 32612 4519 32668
rect 4455 32608 4519 32612
rect 7479 32668 7543 32672
rect 7479 32612 7483 32668
rect 7483 32612 7539 32668
rect 7539 32612 7543 32668
rect 7479 32608 7543 32612
rect 7559 32668 7623 32672
rect 7559 32612 7563 32668
rect 7563 32612 7619 32668
rect 7619 32612 7623 32668
rect 7559 32608 7623 32612
rect 7639 32668 7703 32672
rect 7639 32612 7643 32668
rect 7643 32612 7699 32668
rect 7699 32612 7703 32668
rect 7639 32608 7703 32612
rect 7719 32668 7783 32672
rect 7719 32612 7723 32668
rect 7723 32612 7779 32668
rect 7779 32612 7783 32668
rect 7719 32608 7783 32612
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 5847 32124 5911 32128
rect 5847 32068 5851 32124
rect 5851 32068 5907 32124
rect 5907 32068 5911 32124
rect 5847 32064 5911 32068
rect 5927 32124 5991 32128
rect 5927 32068 5931 32124
rect 5931 32068 5987 32124
rect 5987 32068 5991 32124
rect 5927 32064 5991 32068
rect 6007 32124 6071 32128
rect 6007 32068 6011 32124
rect 6011 32068 6067 32124
rect 6067 32068 6071 32124
rect 6007 32064 6071 32068
rect 6087 32124 6151 32128
rect 6087 32068 6091 32124
rect 6091 32068 6147 32124
rect 6147 32068 6151 32124
rect 6087 32064 6151 32068
rect 9111 32124 9175 32128
rect 9111 32068 9115 32124
rect 9115 32068 9171 32124
rect 9171 32068 9175 32124
rect 9111 32064 9175 32068
rect 9191 32124 9255 32128
rect 9191 32068 9195 32124
rect 9195 32068 9251 32124
rect 9251 32068 9255 32124
rect 9191 32064 9255 32068
rect 9271 32124 9335 32128
rect 9271 32068 9275 32124
rect 9275 32068 9331 32124
rect 9331 32068 9335 32124
rect 9271 32064 9335 32068
rect 9351 32124 9415 32128
rect 9351 32068 9355 32124
rect 9355 32068 9411 32124
rect 9411 32068 9415 32124
rect 9351 32064 9415 32068
rect 3004 31996 3068 32060
rect 1900 31920 1964 31924
rect 1900 31864 1914 31920
rect 1914 31864 1964 31920
rect 1900 31860 1964 31864
rect 2268 31724 2332 31788
rect 4215 31580 4279 31584
rect 4215 31524 4219 31580
rect 4219 31524 4275 31580
rect 4275 31524 4279 31580
rect 4215 31520 4279 31524
rect 4295 31580 4359 31584
rect 4295 31524 4299 31580
rect 4299 31524 4355 31580
rect 4355 31524 4359 31580
rect 4295 31520 4359 31524
rect 4375 31580 4439 31584
rect 4375 31524 4379 31580
rect 4379 31524 4435 31580
rect 4435 31524 4439 31580
rect 4375 31520 4439 31524
rect 4455 31580 4519 31584
rect 4455 31524 4459 31580
rect 4459 31524 4515 31580
rect 4515 31524 4519 31580
rect 4455 31520 4519 31524
rect 7479 31580 7543 31584
rect 7479 31524 7483 31580
rect 7483 31524 7539 31580
rect 7539 31524 7543 31580
rect 7479 31520 7543 31524
rect 7559 31580 7623 31584
rect 7559 31524 7563 31580
rect 7563 31524 7619 31580
rect 7619 31524 7623 31580
rect 7559 31520 7623 31524
rect 7639 31580 7703 31584
rect 7639 31524 7643 31580
rect 7643 31524 7699 31580
rect 7699 31524 7703 31580
rect 7639 31520 7703 31524
rect 7719 31580 7783 31584
rect 7719 31524 7723 31580
rect 7723 31524 7779 31580
rect 7779 31524 7783 31580
rect 7719 31520 7783 31524
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5847 31036 5911 31040
rect 5847 30980 5851 31036
rect 5851 30980 5907 31036
rect 5907 30980 5911 31036
rect 5847 30976 5911 30980
rect 5927 31036 5991 31040
rect 5927 30980 5931 31036
rect 5931 30980 5987 31036
rect 5987 30980 5991 31036
rect 5927 30976 5991 30980
rect 6007 31036 6071 31040
rect 6007 30980 6011 31036
rect 6011 30980 6067 31036
rect 6067 30980 6071 31036
rect 6007 30976 6071 30980
rect 6087 31036 6151 31040
rect 6087 30980 6091 31036
rect 6091 30980 6147 31036
rect 6147 30980 6151 31036
rect 6087 30976 6151 30980
rect 9111 31036 9175 31040
rect 9111 30980 9115 31036
rect 9115 30980 9171 31036
rect 9171 30980 9175 31036
rect 9111 30976 9175 30980
rect 9191 31036 9255 31040
rect 9191 30980 9195 31036
rect 9195 30980 9251 31036
rect 9251 30980 9255 31036
rect 9191 30976 9255 30980
rect 9271 31036 9335 31040
rect 9271 30980 9275 31036
rect 9275 30980 9331 31036
rect 9331 30980 9335 31036
rect 9271 30976 9335 30980
rect 9351 31036 9415 31040
rect 9351 30980 9355 31036
rect 9355 30980 9411 31036
rect 9411 30980 9415 31036
rect 9351 30976 9415 30980
rect 4215 30492 4279 30496
rect 4215 30436 4219 30492
rect 4219 30436 4275 30492
rect 4275 30436 4279 30492
rect 4215 30432 4279 30436
rect 4295 30492 4359 30496
rect 4295 30436 4299 30492
rect 4299 30436 4355 30492
rect 4355 30436 4359 30492
rect 4295 30432 4359 30436
rect 4375 30492 4439 30496
rect 4375 30436 4379 30492
rect 4379 30436 4435 30492
rect 4435 30436 4439 30492
rect 4375 30432 4439 30436
rect 4455 30492 4519 30496
rect 4455 30436 4459 30492
rect 4459 30436 4515 30492
rect 4515 30436 4519 30492
rect 4455 30432 4519 30436
rect 7479 30492 7543 30496
rect 7479 30436 7483 30492
rect 7483 30436 7539 30492
rect 7539 30436 7543 30492
rect 7479 30432 7543 30436
rect 7559 30492 7623 30496
rect 7559 30436 7563 30492
rect 7563 30436 7619 30492
rect 7619 30436 7623 30492
rect 7559 30432 7623 30436
rect 7639 30492 7703 30496
rect 7639 30436 7643 30492
rect 7643 30436 7699 30492
rect 7699 30436 7703 30492
rect 7639 30432 7703 30436
rect 7719 30492 7783 30496
rect 7719 30436 7723 30492
rect 7723 30436 7779 30492
rect 7779 30436 7783 30492
rect 7719 30432 7783 30436
rect 3740 30152 3804 30156
rect 3740 30096 3790 30152
rect 3790 30096 3804 30152
rect 3740 30092 3804 30096
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5847 29948 5911 29952
rect 5847 29892 5851 29948
rect 5851 29892 5907 29948
rect 5907 29892 5911 29948
rect 5847 29888 5911 29892
rect 5927 29948 5991 29952
rect 5927 29892 5931 29948
rect 5931 29892 5987 29948
rect 5987 29892 5991 29948
rect 5927 29888 5991 29892
rect 6007 29948 6071 29952
rect 6007 29892 6011 29948
rect 6011 29892 6067 29948
rect 6067 29892 6071 29948
rect 6007 29888 6071 29892
rect 6087 29948 6151 29952
rect 6087 29892 6091 29948
rect 6091 29892 6147 29948
rect 6147 29892 6151 29948
rect 6087 29888 6151 29892
rect 9111 29948 9175 29952
rect 9111 29892 9115 29948
rect 9115 29892 9171 29948
rect 9171 29892 9175 29948
rect 9111 29888 9175 29892
rect 9191 29948 9255 29952
rect 9191 29892 9195 29948
rect 9195 29892 9251 29948
rect 9251 29892 9255 29948
rect 9191 29888 9255 29892
rect 9271 29948 9335 29952
rect 9271 29892 9275 29948
rect 9275 29892 9331 29948
rect 9331 29892 9335 29948
rect 9271 29888 9335 29892
rect 9351 29948 9415 29952
rect 9351 29892 9355 29948
rect 9355 29892 9411 29948
rect 9411 29892 9415 29948
rect 9351 29888 9415 29892
rect 4215 29404 4279 29408
rect 4215 29348 4219 29404
rect 4219 29348 4275 29404
rect 4275 29348 4279 29404
rect 4215 29344 4279 29348
rect 4295 29404 4359 29408
rect 4295 29348 4299 29404
rect 4299 29348 4355 29404
rect 4355 29348 4359 29404
rect 4295 29344 4359 29348
rect 4375 29404 4439 29408
rect 4375 29348 4379 29404
rect 4379 29348 4435 29404
rect 4435 29348 4439 29404
rect 4375 29344 4439 29348
rect 4455 29404 4519 29408
rect 4455 29348 4459 29404
rect 4459 29348 4515 29404
rect 4515 29348 4519 29404
rect 4455 29344 4519 29348
rect 7479 29404 7543 29408
rect 7479 29348 7483 29404
rect 7483 29348 7539 29404
rect 7539 29348 7543 29404
rect 7479 29344 7543 29348
rect 7559 29404 7623 29408
rect 7559 29348 7563 29404
rect 7563 29348 7619 29404
rect 7619 29348 7623 29404
rect 7559 29344 7623 29348
rect 7639 29404 7703 29408
rect 7639 29348 7643 29404
rect 7643 29348 7699 29404
rect 7699 29348 7703 29404
rect 7639 29344 7703 29348
rect 7719 29404 7783 29408
rect 7719 29348 7723 29404
rect 7723 29348 7779 29404
rect 7779 29348 7783 29404
rect 7719 29344 7783 29348
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5847 28860 5911 28864
rect 5847 28804 5851 28860
rect 5851 28804 5907 28860
rect 5907 28804 5911 28860
rect 5847 28800 5911 28804
rect 5927 28860 5991 28864
rect 5927 28804 5931 28860
rect 5931 28804 5987 28860
rect 5987 28804 5991 28860
rect 5927 28800 5991 28804
rect 6007 28860 6071 28864
rect 6007 28804 6011 28860
rect 6011 28804 6067 28860
rect 6067 28804 6071 28860
rect 6007 28800 6071 28804
rect 6087 28860 6151 28864
rect 6087 28804 6091 28860
rect 6091 28804 6147 28860
rect 6147 28804 6151 28860
rect 6087 28800 6151 28804
rect 9111 28860 9175 28864
rect 9111 28804 9115 28860
rect 9115 28804 9171 28860
rect 9171 28804 9175 28860
rect 9111 28800 9175 28804
rect 9191 28860 9255 28864
rect 9191 28804 9195 28860
rect 9195 28804 9251 28860
rect 9251 28804 9255 28860
rect 9191 28800 9255 28804
rect 9271 28860 9335 28864
rect 9271 28804 9275 28860
rect 9275 28804 9331 28860
rect 9331 28804 9335 28860
rect 9271 28800 9335 28804
rect 9351 28860 9415 28864
rect 9351 28804 9355 28860
rect 9355 28804 9411 28860
rect 9411 28804 9415 28860
rect 9351 28800 9415 28804
rect 3188 28792 3252 28796
rect 3188 28736 3202 28792
rect 3202 28736 3252 28792
rect 3188 28732 3252 28736
rect 4215 28316 4279 28320
rect 4215 28260 4219 28316
rect 4219 28260 4275 28316
rect 4275 28260 4279 28316
rect 4215 28256 4279 28260
rect 4295 28316 4359 28320
rect 4295 28260 4299 28316
rect 4299 28260 4355 28316
rect 4355 28260 4359 28316
rect 4295 28256 4359 28260
rect 4375 28316 4439 28320
rect 4375 28260 4379 28316
rect 4379 28260 4435 28316
rect 4435 28260 4439 28316
rect 4375 28256 4439 28260
rect 4455 28316 4519 28320
rect 4455 28260 4459 28316
rect 4459 28260 4515 28316
rect 4515 28260 4519 28316
rect 4455 28256 4519 28260
rect 7479 28316 7543 28320
rect 7479 28260 7483 28316
rect 7483 28260 7539 28316
rect 7539 28260 7543 28316
rect 7479 28256 7543 28260
rect 7559 28316 7623 28320
rect 7559 28260 7563 28316
rect 7563 28260 7619 28316
rect 7619 28260 7623 28316
rect 7559 28256 7623 28260
rect 7639 28316 7703 28320
rect 7639 28260 7643 28316
rect 7643 28260 7699 28316
rect 7699 28260 7703 28316
rect 7639 28256 7703 28260
rect 7719 28316 7783 28320
rect 7719 28260 7723 28316
rect 7723 28260 7779 28316
rect 7779 28260 7783 28316
rect 7719 28256 7783 28260
rect 1900 28052 1964 28116
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5847 27772 5911 27776
rect 5847 27716 5851 27772
rect 5851 27716 5907 27772
rect 5907 27716 5911 27772
rect 5847 27712 5911 27716
rect 5927 27772 5991 27776
rect 5927 27716 5931 27772
rect 5931 27716 5987 27772
rect 5987 27716 5991 27772
rect 5927 27712 5991 27716
rect 6007 27772 6071 27776
rect 6007 27716 6011 27772
rect 6011 27716 6067 27772
rect 6067 27716 6071 27772
rect 6007 27712 6071 27716
rect 6087 27772 6151 27776
rect 6087 27716 6091 27772
rect 6091 27716 6147 27772
rect 6147 27716 6151 27772
rect 6087 27712 6151 27716
rect 9111 27772 9175 27776
rect 9111 27716 9115 27772
rect 9115 27716 9171 27772
rect 9171 27716 9175 27772
rect 9111 27712 9175 27716
rect 9191 27772 9255 27776
rect 9191 27716 9195 27772
rect 9195 27716 9251 27772
rect 9251 27716 9255 27772
rect 9191 27712 9255 27716
rect 9271 27772 9335 27776
rect 9271 27716 9275 27772
rect 9275 27716 9331 27772
rect 9331 27716 9335 27772
rect 9271 27712 9335 27716
rect 9351 27772 9415 27776
rect 9351 27716 9355 27772
rect 9355 27716 9411 27772
rect 9411 27716 9415 27772
rect 9351 27712 9415 27716
rect 3004 27508 3068 27572
rect 4215 27228 4279 27232
rect 4215 27172 4219 27228
rect 4219 27172 4275 27228
rect 4275 27172 4279 27228
rect 4215 27168 4279 27172
rect 4295 27228 4359 27232
rect 4295 27172 4299 27228
rect 4299 27172 4355 27228
rect 4355 27172 4359 27228
rect 4295 27168 4359 27172
rect 4375 27228 4439 27232
rect 4375 27172 4379 27228
rect 4379 27172 4435 27228
rect 4435 27172 4439 27228
rect 4375 27168 4439 27172
rect 4455 27228 4519 27232
rect 4455 27172 4459 27228
rect 4459 27172 4515 27228
rect 4515 27172 4519 27228
rect 4455 27168 4519 27172
rect 7479 27228 7543 27232
rect 7479 27172 7483 27228
rect 7483 27172 7539 27228
rect 7539 27172 7543 27228
rect 7479 27168 7543 27172
rect 7559 27228 7623 27232
rect 7559 27172 7563 27228
rect 7563 27172 7619 27228
rect 7619 27172 7623 27228
rect 7559 27168 7623 27172
rect 7639 27228 7703 27232
rect 7639 27172 7643 27228
rect 7643 27172 7699 27228
rect 7699 27172 7703 27228
rect 7639 27168 7703 27172
rect 7719 27228 7783 27232
rect 7719 27172 7723 27228
rect 7723 27172 7779 27228
rect 7779 27172 7783 27228
rect 7719 27168 7783 27172
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5847 26684 5911 26688
rect 5847 26628 5851 26684
rect 5851 26628 5907 26684
rect 5907 26628 5911 26684
rect 5847 26624 5911 26628
rect 5927 26684 5991 26688
rect 5927 26628 5931 26684
rect 5931 26628 5987 26684
rect 5987 26628 5991 26684
rect 5927 26624 5991 26628
rect 6007 26684 6071 26688
rect 6007 26628 6011 26684
rect 6011 26628 6067 26684
rect 6067 26628 6071 26684
rect 6007 26624 6071 26628
rect 6087 26684 6151 26688
rect 6087 26628 6091 26684
rect 6091 26628 6147 26684
rect 6147 26628 6151 26684
rect 6087 26624 6151 26628
rect 9111 26684 9175 26688
rect 9111 26628 9115 26684
rect 9115 26628 9171 26684
rect 9171 26628 9175 26684
rect 9111 26624 9175 26628
rect 9191 26684 9255 26688
rect 9191 26628 9195 26684
rect 9195 26628 9251 26684
rect 9251 26628 9255 26684
rect 9191 26624 9255 26628
rect 9271 26684 9335 26688
rect 9271 26628 9275 26684
rect 9275 26628 9331 26684
rect 9331 26628 9335 26684
rect 9271 26624 9335 26628
rect 9351 26684 9415 26688
rect 9351 26628 9355 26684
rect 9355 26628 9411 26684
rect 9411 26628 9415 26684
rect 9351 26624 9415 26628
rect 4215 26140 4279 26144
rect 4215 26084 4219 26140
rect 4219 26084 4275 26140
rect 4275 26084 4279 26140
rect 4215 26080 4279 26084
rect 4295 26140 4359 26144
rect 4295 26084 4299 26140
rect 4299 26084 4355 26140
rect 4355 26084 4359 26140
rect 4295 26080 4359 26084
rect 4375 26140 4439 26144
rect 4375 26084 4379 26140
rect 4379 26084 4435 26140
rect 4435 26084 4439 26140
rect 4375 26080 4439 26084
rect 4455 26140 4519 26144
rect 4455 26084 4459 26140
rect 4459 26084 4515 26140
rect 4515 26084 4519 26140
rect 4455 26080 4519 26084
rect 7479 26140 7543 26144
rect 7479 26084 7483 26140
rect 7483 26084 7539 26140
rect 7539 26084 7543 26140
rect 7479 26080 7543 26084
rect 7559 26140 7623 26144
rect 7559 26084 7563 26140
rect 7563 26084 7619 26140
rect 7619 26084 7623 26140
rect 7559 26080 7623 26084
rect 7639 26140 7703 26144
rect 7639 26084 7643 26140
rect 7643 26084 7699 26140
rect 7699 26084 7703 26140
rect 7639 26080 7703 26084
rect 7719 26140 7783 26144
rect 7719 26084 7723 26140
rect 7723 26084 7779 26140
rect 7779 26084 7783 26140
rect 7719 26080 7783 26084
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5847 25596 5911 25600
rect 5847 25540 5851 25596
rect 5851 25540 5907 25596
rect 5907 25540 5911 25596
rect 5847 25536 5911 25540
rect 5927 25596 5991 25600
rect 5927 25540 5931 25596
rect 5931 25540 5987 25596
rect 5987 25540 5991 25596
rect 5927 25536 5991 25540
rect 6007 25596 6071 25600
rect 6007 25540 6011 25596
rect 6011 25540 6067 25596
rect 6067 25540 6071 25596
rect 6007 25536 6071 25540
rect 6087 25596 6151 25600
rect 6087 25540 6091 25596
rect 6091 25540 6147 25596
rect 6147 25540 6151 25596
rect 6087 25536 6151 25540
rect 9111 25596 9175 25600
rect 9111 25540 9115 25596
rect 9115 25540 9171 25596
rect 9171 25540 9175 25596
rect 9111 25536 9175 25540
rect 9191 25596 9255 25600
rect 9191 25540 9195 25596
rect 9195 25540 9251 25596
rect 9251 25540 9255 25596
rect 9191 25536 9255 25540
rect 9271 25596 9335 25600
rect 9271 25540 9275 25596
rect 9275 25540 9331 25596
rect 9331 25540 9335 25596
rect 9271 25536 9335 25540
rect 9351 25596 9415 25600
rect 9351 25540 9355 25596
rect 9355 25540 9411 25596
rect 9411 25540 9415 25596
rect 9351 25536 9415 25540
rect 4215 25052 4279 25056
rect 4215 24996 4219 25052
rect 4219 24996 4275 25052
rect 4275 24996 4279 25052
rect 4215 24992 4279 24996
rect 4295 25052 4359 25056
rect 4295 24996 4299 25052
rect 4299 24996 4355 25052
rect 4355 24996 4359 25052
rect 4295 24992 4359 24996
rect 4375 25052 4439 25056
rect 4375 24996 4379 25052
rect 4379 24996 4435 25052
rect 4435 24996 4439 25052
rect 4375 24992 4439 24996
rect 4455 25052 4519 25056
rect 4455 24996 4459 25052
rect 4459 24996 4515 25052
rect 4515 24996 4519 25052
rect 4455 24992 4519 24996
rect 7479 25052 7543 25056
rect 7479 24996 7483 25052
rect 7483 24996 7539 25052
rect 7539 24996 7543 25052
rect 7479 24992 7543 24996
rect 7559 25052 7623 25056
rect 7559 24996 7563 25052
rect 7563 24996 7619 25052
rect 7619 24996 7623 25052
rect 7559 24992 7623 24996
rect 7639 25052 7703 25056
rect 7639 24996 7643 25052
rect 7643 24996 7699 25052
rect 7699 24996 7703 25052
rect 7639 24992 7703 24996
rect 7719 25052 7783 25056
rect 7719 24996 7723 25052
rect 7723 24996 7779 25052
rect 7779 24996 7783 25052
rect 7719 24992 7783 24996
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5847 24508 5911 24512
rect 5847 24452 5851 24508
rect 5851 24452 5907 24508
rect 5907 24452 5911 24508
rect 5847 24448 5911 24452
rect 5927 24508 5991 24512
rect 5927 24452 5931 24508
rect 5931 24452 5987 24508
rect 5987 24452 5991 24508
rect 5927 24448 5991 24452
rect 6007 24508 6071 24512
rect 6007 24452 6011 24508
rect 6011 24452 6067 24508
rect 6067 24452 6071 24508
rect 6007 24448 6071 24452
rect 6087 24508 6151 24512
rect 6087 24452 6091 24508
rect 6091 24452 6147 24508
rect 6147 24452 6151 24508
rect 6087 24448 6151 24452
rect 9111 24508 9175 24512
rect 9111 24452 9115 24508
rect 9115 24452 9171 24508
rect 9171 24452 9175 24508
rect 9111 24448 9175 24452
rect 9191 24508 9255 24512
rect 9191 24452 9195 24508
rect 9195 24452 9251 24508
rect 9251 24452 9255 24508
rect 9191 24448 9255 24452
rect 9271 24508 9335 24512
rect 9271 24452 9275 24508
rect 9275 24452 9331 24508
rect 9331 24452 9335 24508
rect 9271 24448 9335 24452
rect 9351 24508 9415 24512
rect 9351 24452 9355 24508
rect 9355 24452 9411 24508
rect 9411 24452 9415 24508
rect 9351 24448 9415 24452
rect 4215 23964 4279 23968
rect 4215 23908 4219 23964
rect 4219 23908 4275 23964
rect 4275 23908 4279 23964
rect 4215 23904 4279 23908
rect 4295 23964 4359 23968
rect 4295 23908 4299 23964
rect 4299 23908 4355 23964
rect 4355 23908 4359 23964
rect 4295 23904 4359 23908
rect 4375 23964 4439 23968
rect 4375 23908 4379 23964
rect 4379 23908 4435 23964
rect 4435 23908 4439 23964
rect 4375 23904 4439 23908
rect 4455 23964 4519 23968
rect 4455 23908 4459 23964
rect 4459 23908 4515 23964
rect 4515 23908 4519 23964
rect 4455 23904 4519 23908
rect 7479 23964 7543 23968
rect 7479 23908 7483 23964
rect 7483 23908 7539 23964
rect 7539 23908 7543 23964
rect 7479 23904 7543 23908
rect 7559 23964 7623 23968
rect 7559 23908 7563 23964
rect 7563 23908 7619 23964
rect 7619 23908 7623 23964
rect 7559 23904 7623 23908
rect 7639 23964 7703 23968
rect 7639 23908 7643 23964
rect 7643 23908 7699 23964
rect 7699 23908 7703 23964
rect 7639 23904 7703 23908
rect 7719 23964 7783 23968
rect 7719 23908 7723 23964
rect 7723 23908 7779 23964
rect 7779 23908 7783 23964
rect 7719 23904 7783 23908
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5847 23420 5911 23424
rect 5847 23364 5851 23420
rect 5851 23364 5907 23420
rect 5907 23364 5911 23420
rect 5847 23360 5911 23364
rect 5927 23420 5991 23424
rect 5927 23364 5931 23420
rect 5931 23364 5987 23420
rect 5987 23364 5991 23420
rect 5927 23360 5991 23364
rect 6007 23420 6071 23424
rect 6007 23364 6011 23420
rect 6011 23364 6067 23420
rect 6067 23364 6071 23420
rect 6007 23360 6071 23364
rect 6087 23420 6151 23424
rect 6087 23364 6091 23420
rect 6091 23364 6147 23420
rect 6147 23364 6151 23420
rect 6087 23360 6151 23364
rect 9111 23420 9175 23424
rect 9111 23364 9115 23420
rect 9115 23364 9171 23420
rect 9171 23364 9175 23420
rect 9111 23360 9175 23364
rect 9191 23420 9255 23424
rect 9191 23364 9195 23420
rect 9195 23364 9251 23420
rect 9251 23364 9255 23420
rect 9191 23360 9255 23364
rect 9271 23420 9335 23424
rect 9271 23364 9275 23420
rect 9275 23364 9331 23420
rect 9331 23364 9335 23420
rect 9271 23360 9335 23364
rect 9351 23420 9415 23424
rect 9351 23364 9355 23420
rect 9355 23364 9411 23420
rect 9411 23364 9415 23420
rect 9351 23360 9415 23364
rect 4215 22876 4279 22880
rect 4215 22820 4219 22876
rect 4219 22820 4275 22876
rect 4275 22820 4279 22876
rect 4215 22816 4279 22820
rect 4295 22876 4359 22880
rect 4295 22820 4299 22876
rect 4299 22820 4355 22876
rect 4355 22820 4359 22876
rect 4295 22816 4359 22820
rect 4375 22876 4439 22880
rect 4375 22820 4379 22876
rect 4379 22820 4435 22876
rect 4435 22820 4439 22876
rect 4375 22816 4439 22820
rect 4455 22876 4519 22880
rect 4455 22820 4459 22876
rect 4459 22820 4515 22876
rect 4515 22820 4519 22876
rect 4455 22816 4519 22820
rect 7479 22876 7543 22880
rect 7479 22820 7483 22876
rect 7483 22820 7539 22876
rect 7539 22820 7543 22876
rect 7479 22816 7543 22820
rect 7559 22876 7623 22880
rect 7559 22820 7563 22876
rect 7563 22820 7619 22876
rect 7619 22820 7623 22876
rect 7559 22816 7623 22820
rect 7639 22876 7703 22880
rect 7639 22820 7643 22876
rect 7643 22820 7699 22876
rect 7699 22820 7703 22876
rect 7639 22816 7703 22820
rect 7719 22876 7783 22880
rect 7719 22820 7723 22876
rect 7723 22820 7779 22876
rect 7779 22820 7783 22876
rect 7719 22816 7783 22820
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5847 22332 5911 22336
rect 5847 22276 5851 22332
rect 5851 22276 5907 22332
rect 5907 22276 5911 22332
rect 5847 22272 5911 22276
rect 5927 22332 5991 22336
rect 5927 22276 5931 22332
rect 5931 22276 5987 22332
rect 5987 22276 5991 22332
rect 5927 22272 5991 22276
rect 6007 22332 6071 22336
rect 6007 22276 6011 22332
rect 6011 22276 6067 22332
rect 6067 22276 6071 22332
rect 6007 22272 6071 22276
rect 6087 22332 6151 22336
rect 6087 22276 6091 22332
rect 6091 22276 6147 22332
rect 6147 22276 6151 22332
rect 6087 22272 6151 22276
rect 9111 22332 9175 22336
rect 9111 22276 9115 22332
rect 9115 22276 9171 22332
rect 9171 22276 9175 22332
rect 9111 22272 9175 22276
rect 9191 22332 9255 22336
rect 9191 22276 9195 22332
rect 9195 22276 9251 22332
rect 9251 22276 9255 22332
rect 9191 22272 9255 22276
rect 9271 22332 9335 22336
rect 9271 22276 9275 22332
rect 9275 22276 9331 22332
rect 9331 22276 9335 22332
rect 9271 22272 9335 22276
rect 9351 22332 9415 22336
rect 9351 22276 9355 22332
rect 9355 22276 9411 22332
rect 9411 22276 9415 22332
rect 9351 22272 9415 22276
rect 3188 21932 3252 21996
rect 4215 21788 4279 21792
rect 4215 21732 4219 21788
rect 4219 21732 4275 21788
rect 4275 21732 4279 21788
rect 4215 21728 4279 21732
rect 4295 21788 4359 21792
rect 4295 21732 4299 21788
rect 4299 21732 4355 21788
rect 4355 21732 4359 21788
rect 4295 21728 4359 21732
rect 4375 21788 4439 21792
rect 4375 21732 4379 21788
rect 4379 21732 4435 21788
rect 4435 21732 4439 21788
rect 4375 21728 4439 21732
rect 4455 21788 4519 21792
rect 4455 21732 4459 21788
rect 4459 21732 4515 21788
rect 4515 21732 4519 21788
rect 4455 21728 4519 21732
rect 7479 21788 7543 21792
rect 7479 21732 7483 21788
rect 7483 21732 7539 21788
rect 7539 21732 7543 21788
rect 7479 21728 7543 21732
rect 7559 21788 7623 21792
rect 7559 21732 7563 21788
rect 7563 21732 7619 21788
rect 7619 21732 7623 21788
rect 7559 21728 7623 21732
rect 7639 21788 7703 21792
rect 7639 21732 7643 21788
rect 7643 21732 7699 21788
rect 7699 21732 7703 21788
rect 7639 21728 7703 21732
rect 7719 21788 7783 21792
rect 7719 21732 7723 21788
rect 7723 21732 7779 21788
rect 7779 21732 7783 21788
rect 7719 21728 7783 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5847 21244 5911 21248
rect 5847 21188 5851 21244
rect 5851 21188 5907 21244
rect 5907 21188 5911 21244
rect 5847 21184 5911 21188
rect 5927 21244 5991 21248
rect 5927 21188 5931 21244
rect 5931 21188 5987 21244
rect 5987 21188 5991 21244
rect 5927 21184 5991 21188
rect 6007 21244 6071 21248
rect 6007 21188 6011 21244
rect 6011 21188 6067 21244
rect 6067 21188 6071 21244
rect 6007 21184 6071 21188
rect 6087 21244 6151 21248
rect 6087 21188 6091 21244
rect 6091 21188 6147 21244
rect 6147 21188 6151 21244
rect 6087 21184 6151 21188
rect 9111 21244 9175 21248
rect 9111 21188 9115 21244
rect 9115 21188 9171 21244
rect 9171 21188 9175 21244
rect 9111 21184 9175 21188
rect 9191 21244 9255 21248
rect 9191 21188 9195 21244
rect 9195 21188 9251 21244
rect 9251 21188 9255 21244
rect 9191 21184 9255 21188
rect 9271 21244 9335 21248
rect 9271 21188 9275 21244
rect 9275 21188 9331 21244
rect 9331 21188 9335 21244
rect 9271 21184 9335 21188
rect 9351 21244 9415 21248
rect 9351 21188 9355 21244
rect 9355 21188 9411 21244
rect 9411 21188 9415 21244
rect 9351 21184 9415 21188
rect 4215 20700 4279 20704
rect 4215 20644 4219 20700
rect 4219 20644 4275 20700
rect 4275 20644 4279 20700
rect 4215 20640 4279 20644
rect 4295 20700 4359 20704
rect 4295 20644 4299 20700
rect 4299 20644 4355 20700
rect 4355 20644 4359 20700
rect 4295 20640 4359 20644
rect 4375 20700 4439 20704
rect 4375 20644 4379 20700
rect 4379 20644 4435 20700
rect 4435 20644 4439 20700
rect 4375 20640 4439 20644
rect 4455 20700 4519 20704
rect 4455 20644 4459 20700
rect 4459 20644 4515 20700
rect 4515 20644 4519 20700
rect 4455 20640 4519 20644
rect 7479 20700 7543 20704
rect 7479 20644 7483 20700
rect 7483 20644 7539 20700
rect 7539 20644 7543 20700
rect 7479 20640 7543 20644
rect 7559 20700 7623 20704
rect 7559 20644 7563 20700
rect 7563 20644 7619 20700
rect 7619 20644 7623 20700
rect 7559 20640 7623 20644
rect 7639 20700 7703 20704
rect 7639 20644 7643 20700
rect 7643 20644 7699 20700
rect 7699 20644 7703 20700
rect 7639 20640 7703 20644
rect 7719 20700 7783 20704
rect 7719 20644 7723 20700
rect 7723 20644 7779 20700
rect 7779 20644 7783 20700
rect 7719 20640 7783 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5847 20156 5911 20160
rect 5847 20100 5851 20156
rect 5851 20100 5907 20156
rect 5907 20100 5911 20156
rect 5847 20096 5911 20100
rect 5927 20156 5991 20160
rect 5927 20100 5931 20156
rect 5931 20100 5987 20156
rect 5987 20100 5991 20156
rect 5927 20096 5991 20100
rect 6007 20156 6071 20160
rect 6007 20100 6011 20156
rect 6011 20100 6067 20156
rect 6067 20100 6071 20156
rect 6007 20096 6071 20100
rect 6087 20156 6151 20160
rect 6087 20100 6091 20156
rect 6091 20100 6147 20156
rect 6147 20100 6151 20156
rect 6087 20096 6151 20100
rect 9111 20156 9175 20160
rect 9111 20100 9115 20156
rect 9115 20100 9171 20156
rect 9171 20100 9175 20156
rect 9111 20096 9175 20100
rect 9191 20156 9255 20160
rect 9191 20100 9195 20156
rect 9195 20100 9251 20156
rect 9251 20100 9255 20156
rect 9191 20096 9255 20100
rect 9271 20156 9335 20160
rect 9271 20100 9275 20156
rect 9275 20100 9331 20156
rect 9331 20100 9335 20156
rect 9271 20096 9335 20100
rect 9351 20156 9415 20160
rect 9351 20100 9355 20156
rect 9355 20100 9411 20156
rect 9411 20100 9415 20156
rect 9351 20096 9415 20100
rect 4215 19612 4279 19616
rect 4215 19556 4219 19612
rect 4219 19556 4275 19612
rect 4275 19556 4279 19612
rect 4215 19552 4279 19556
rect 4295 19612 4359 19616
rect 4295 19556 4299 19612
rect 4299 19556 4355 19612
rect 4355 19556 4359 19612
rect 4295 19552 4359 19556
rect 4375 19612 4439 19616
rect 4375 19556 4379 19612
rect 4379 19556 4435 19612
rect 4435 19556 4439 19612
rect 4375 19552 4439 19556
rect 4455 19612 4519 19616
rect 4455 19556 4459 19612
rect 4459 19556 4515 19612
rect 4515 19556 4519 19612
rect 4455 19552 4519 19556
rect 7479 19612 7543 19616
rect 7479 19556 7483 19612
rect 7483 19556 7539 19612
rect 7539 19556 7543 19612
rect 7479 19552 7543 19556
rect 7559 19612 7623 19616
rect 7559 19556 7563 19612
rect 7563 19556 7619 19612
rect 7619 19556 7623 19612
rect 7559 19552 7623 19556
rect 7639 19612 7703 19616
rect 7639 19556 7643 19612
rect 7643 19556 7699 19612
rect 7699 19556 7703 19612
rect 7639 19552 7703 19556
rect 7719 19612 7783 19616
rect 7719 19556 7723 19612
rect 7723 19556 7779 19612
rect 7779 19556 7783 19612
rect 7719 19552 7783 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5847 19068 5911 19072
rect 5847 19012 5851 19068
rect 5851 19012 5907 19068
rect 5907 19012 5911 19068
rect 5847 19008 5911 19012
rect 5927 19068 5991 19072
rect 5927 19012 5931 19068
rect 5931 19012 5987 19068
rect 5987 19012 5991 19068
rect 5927 19008 5991 19012
rect 6007 19068 6071 19072
rect 6007 19012 6011 19068
rect 6011 19012 6067 19068
rect 6067 19012 6071 19068
rect 6007 19008 6071 19012
rect 6087 19068 6151 19072
rect 6087 19012 6091 19068
rect 6091 19012 6147 19068
rect 6147 19012 6151 19068
rect 6087 19008 6151 19012
rect 9111 19068 9175 19072
rect 9111 19012 9115 19068
rect 9115 19012 9171 19068
rect 9171 19012 9175 19068
rect 9111 19008 9175 19012
rect 9191 19068 9255 19072
rect 9191 19012 9195 19068
rect 9195 19012 9251 19068
rect 9251 19012 9255 19068
rect 9191 19008 9255 19012
rect 9271 19068 9335 19072
rect 9271 19012 9275 19068
rect 9275 19012 9331 19068
rect 9331 19012 9335 19068
rect 9271 19008 9335 19012
rect 9351 19068 9415 19072
rect 9351 19012 9355 19068
rect 9355 19012 9411 19068
rect 9411 19012 9415 19068
rect 9351 19008 9415 19012
rect 4215 18524 4279 18528
rect 4215 18468 4219 18524
rect 4219 18468 4275 18524
rect 4275 18468 4279 18524
rect 4215 18464 4279 18468
rect 4295 18524 4359 18528
rect 4295 18468 4299 18524
rect 4299 18468 4355 18524
rect 4355 18468 4359 18524
rect 4295 18464 4359 18468
rect 4375 18524 4439 18528
rect 4375 18468 4379 18524
rect 4379 18468 4435 18524
rect 4435 18468 4439 18524
rect 4375 18464 4439 18468
rect 4455 18524 4519 18528
rect 4455 18468 4459 18524
rect 4459 18468 4515 18524
rect 4515 18468 4519 18524
rect 4455 18464 4519 18468
rect 7479 18524 7543 18528
rect 7479 18468 7483 18524
rect 7483 18468 7539 18524
rect 7539 18468 7543 18524
rect 7479 18464 7543 18468
rect 7559 18524 7623 18528
rect 7559 18468 7563 18524
rect 7563 18468 7619 18524
rect 7619 18468 7623 18524
rect 7559 18464 7623 18468
rect 7639 18524 7703 18528
rect 7639 18468 7643 18524
rect 7643 18468 7699 18524
rect 7699 18468 7703 18524
rect 7639 18464 7703 18468
rect 7719 18524 7783 18528
rect 7719 18468 7723 18524
rect 7723 18468 7779 18524
rect 7779 18468 7783 18524
rect 7719 18464 7783 18468
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5847 17980 5911 17984
rect 5847 17924 5851 17980
rect 5851 17924 5907 17980
rect 5907 17924 5911 17980
rect 5847 17920 5911 17924
rect 5927 17980 5991 17984
rect 5927 17924 5931 17980
rect 5931 17924 5987 17980
rect 5987 17924 5991 17980
rect 5927 17920 5991 17924
rect 6007 17980 6071 17984
rect 6007 17924 6011 17980
rect 6011 17924 6067 17980
rect 6067 17924 6071 17980
rect 6007 17920 6071 17924
rect 6087 17980 6151 17984
rect 6087 17924 6091 17980
rect 6091 17924 6147 17980
rect 6147 17924 6151 17980
rect 6087 17920 6151 17924
rect 9111 17980 9175 17984
rect 9111 17924 9115 17980
rect 9115 17924 9171 17980
rect 9171 17924 9175 17980
rect 9111 17920 9175 17924
rect 9191 17980 9255 17984
rect 9191 17924 9195 17980
rect 9195 17924 9251 17980
rect 9251 17924 9255 17980
rect 9191 17920 9255 17924
rect 9271 17980 9335 17984
rect 9271 17924 9275 17980
rect 9275 17924 9331 17980
rect 9331 17924 9335 17980
rect 9271 17920 9335 17924
rect 9351 17980 9415 17984
rect 9351 17924 9355 17980
rect 9355 17924 9411 17980
rect 9411 17924 9415 17980
rect 9351 17920 9415 17924
rect 4215 17436 4279 17440
rect 4215 17380 4219 17436
rect 4219 17380 4275 17436
rect 4275 17380 4279 17436
rect 4215 17376 4279 17380
rect 4295 17436 4359 17440
rect 4295 17380 4299 17436
rect 4299 17380 4355 17436
rect 4355 17380 4359 17436
rect 4295 17376 4359 17380
rect 4375 17436 4439 17440
rect 4375 17380 4379 17436
rect 4379 17380 4435 17436
rect 4435 17380 4439 17436
rect 4375 17376 4439 17380
rect 4455 17436 4519 17440
rect 4455 17380 4459 17436
rect 4459 17380 4515 17436
rect 4515 17380 4519 17436
rect 4455 17376 4519 17380
rect 7479 17436 7543 17440
rect 7479 17380 7483 17436
rect 7483 17380 7539 17436
rect 7539 17380 7543 17436
rect 7479 17376 7543 17380
rect 7559 17436 7623 17440
rect 7559 17380 7563 17436
rect 7563 17380 7619 17436
rect 7619 17380 7623 17436
rect 7559 17376 7623 17380
rect 7639 17436 7703 17440
rect 7639 17380 7643 17436
rect 7643 17380 7699 17436
rect 7699 17380 7703 17436
rect 7639 17376 7703 17380
rect 7719 17436 7783 17440
rect 7719 17380 7723 17436
rect 7723 17380 7779 17436
rect 7779 17380 7783 17436
rect 7719 17376 7783 17380
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5847 16892 5911 16896
rect 5847 16836 5851 16892
rect 5851 16836 5907 16892
rect 5907 16836 5911 16892
rect 5847 16832 5911 16836
rect 5927 16892 5991 16896
rect 5927 16836 5931 16892
rect 5931 16836 5987 16892
rect 5987 16836 5991 16892
rect 5927 16832 5991 16836
rect 6007 16892 6071 16896
rect 6007 16836 6011 16892
rect 6011 16836 6067 16892
rect 6067 16836 6071 16892
rect 6007 16832 6071 16836
rect 6087 16892 6151 16896
rect 6087 16836 6091 16892
rect 6091 16836 6147 16892
rect 6147 16836 6151 16892
rect 6087 16832 6151 16836
rect 9111 16892 9175 16896
rect 9111 16836 9115 16892
rect 9115 16836 9171 16892
rect 9171 16836 9175 16892
rect 9111 16832 9175 16836
rect 9191 16892 9255 16896
rect 9191 16836 9195 16892
rect 9195 16836 9251 16892
rect 9251 16836 9255 16892
rect 9191 16832 9255 16836
rect 9271 16892 9335 16896
rect 9271 16836 9275 16892
rect 9275 16836 9331 16892
rect 9331 16836 9335 16892
rect 9271 16832 9335 16836
rect 9351 16892 9415 16896
rect 9351 16836 9355 16892
rect 9355 16836 9411 16892
rect 9411 16836 9415 16892
rect 9351 16832 9415 16836
rect 4215 16348 4279 16352
rect 4215 16292 4219 16348
rect 4219 16292 4275 16348
rect 4275 16292 4279 16348
rect 4215 16288 4279 16292
rect 4295 16348 4359 16352
rect 4295 16292 4299 16348
rect 4299 16292 4355 16348
rect 4355 16292 4359 16348
rect 4295 16288 4359 16292
rect 4375 16348 4439 16352
rect 4375 16292 4379 16348
rect 4379 16292 4435 16348
rect 4435 16292 4439 16348
rect 4375 16288 4439 16292
rect 4455 16348 4519 16352
rect 4455 16292 4459 16348
rect 4459 16292 4515 16348
rect 4515 16292 4519 16348
rect 4455 16288 4519 16292
rect 7479 16348 7543 16352
rect 7479 16292 7483 16348
rect 7483 16292 7539 16348
rect 7539 16292 7543 16348
rect 7479 16288 7543 16292
rect 7559 16348 7623 16352
rect 7559 16292 7563 16348
rect 7563 16292 7619 16348
rect 7619 16292 7623 16348
rect 7559 16288 7623 16292
rect 7639 16348 7703 16352
rect 7639 16292 7643 16348
rect 7643 16292 7699 16348
rect 7699 16292 7703 16348
rect 7639 16288 7703 16292
rect 7719 16348 7783 16352
rect 7719 16292 7723 16348
rect 7723 16292 7779 16348
rect 7779 16292 7783 16348
rect 7719 16288 7783 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5847 15804 5911 15808
rect 5847 15748 5851 15804
rect 5851 15748 5907 15804
rect 5907 15748 5911 15804
rect 5847 15744 5911 15748
rect 5927 15804 5991 15808
rect 5927 15748 5931 15804
rect 5931 15748 5987 15804
rect 5987 15748 5991 15804
rect 5927 15744 5991 15748
rect 6007 15804 6071 15808
rect 6007 15748 6011 15804
rect 6011 15748 6067 15804
rect 6067 15748 6071 15804
rect 6007 15744 6071 15748
rect 6087 15804 6151 15808
rect 6087 15748 6091 15804
rect 6091 15748 6147 15804
rect 6147 15748 6151 15804
rect 6087 15744 6151 15748
rect 9111 15804 9175 15808
rect 9111 15748 9115 15804
rect 9115 15748 9171 15804
rect 9171 15748 9175 15804
rect 9111 15744 9175 15748
rect 9191 15804 9255 15808
rect 9191 15748 9195 15804
rect 9195 15748 9251 15804
rect 9251 15748 9255 15804
rect 9191 15744 9255 15748
rect 9271 15804 9335 15808
rect 9271 15748 9275 15804
rect 9275 15748 9331 15804
rect 9331 15748 9335 15804
rect 9271 15744 9335 15748
rect 9351 15804 9415 15808
rect 9351 15748 9355 15804
rect 9355 15748 9411 15804
rect 9411 15748 9415 15804
rect 9351 15744 9415 15748
rect 4215 15260 4279 15264
rect 4215 15204 4219 15260
rect 4219 15204 4275 15260
rect 4275 15204 4279 15260
rect 4215 15200 4279 15204
rect 4295 15260 4359 15264
rect 4295 15204 4299 15260
rect 4299 15204 4355 15260
rect 4355 15204 4359 15260
rect 4295 15200 4359 15204
rect 4375 15260 4439 15264
rect 4375 15204 4379 15260
rect 4379 15204 4435 15260
rect 4435 15204 4439 15260
rect 4375 15200 4439 15204
rect 4455 15260 4519 15264
rect 4455 15204 4459 15260
rect 4459 15204 4515 15260
rect 4515 15204 4519 15260
rect 4455 15200 4519 15204
rect 7479 15260 7543 15264
rect 7479 15204 7483 15260
rect 7483 15204 7539 15260
rect 7539 15204 7543 15260
rect 7479 15200 7543 15204
rect 7559 15260 7623 15264
rect 7559 15204 7563 15260
rect 7563 15204 7619 15260
rect 7619 15204 7623 15260
rect 7559 15200 7623 15204
rect 7639 15260 7703 15264
rect 7639 15204 7643 15260
rect 7643 15204 7699 15260
rect 7699 15204 7703 15260
rect 7639 15200 7703 15204
rect 7719 15260 7783 15264
rect 7719 15204 7723 15260
rect 7723 15204 7779 15260
rect 7779 15204 7783 15260
rect 7719 15200 7783 15204
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5847 14716 5911 14720
rect 5847 14660 5851 14716
rect 5851 14660 5907 14716
rect 5907 14660 5911 14716
rect 5847 14656 5911 14660
rect 5927 14716 5991 14720
rect 5927 14660 5931 14716
rect 5931 14660 5987 14716
rect 5987 14660 5991 14716
rect 5927 14656 5991 14660
rect 6007 14716 6071 14720
rect 6007 14660 6011 14716
rect 6011 14660 6067 14716
rect 6067 14660 6071 14716
rect 6007 14656 6071 14660
rect 6087 14716 6151 14720
rect 6087 14660 6091 14716
rect 6091 14660 6147 14716
rect 6147 14660 6151 14716
rect 6087 14656 6151 14660
rect 9111 14716 9175 14720
rect 9111 14660 9115 14716
rect 9115 14660 9171 14716
rect 9171 14660 9175 14716
rect 9111 14656 9175 14660
rect 9191 14716 9255 14720
rect 9191 14660 9195 14716
rect 9195 14660 9251 14716
rect 9251 14660 9255 14716
rect 9191 14656 9255 14660
rect 9271 14716 9335 14720
rect 9271 14660 9275 14716
rect 9275 14660 9331 14716
rect 9331 14660 9335 14716
rect 9271 14656 9335 14660
rect 9351 14716 9415 14720
rect 9351 14660 9355 14716
rect 9355 14660 9411 14716
rect 9411 14660 9415 14716
rect 9351 14656 9415 14660
rect 4215 14172 4279 14176
rect 4215 14116 4219 14172
rect 4219 14116 4275 14172
rect 4275 14116 4279 14172
rect 4215 14112 4279 14116
rect 4295 14172 4359 14176
rect 4295 14116 4299 14172
rect 4299 14116 4355 14172
rect 4355 14116 4359 14172
rect 4295 14112 4359 14116
rect 4375 14172 4439 14176
rect 4375 14116 4379 14172
rect 4379 14116 4435 14172
rect 4435 14116 4439 14172
rect 4375 14112 4439 14116
rect 4455 14172 4519 14176
rect 4455 14116 4459 14172
rect 4459 14116 4515 14172
rect 4515 14116 4519 14172
rect 4455 14112 4519 14116
rect 7479 14172 7543 14176
rect 7479 14116 7483 14172
rect 7483 14116 7539 14172
rect 7539 14116 7543 14172
rect 7479 14112 7543 14116
rect 7559 14172 7623 14176
rect 7559 14116 7563 14172
rect 7563 14116 7619 14172
rect 7619 14116 7623 14172
rect 7559 14112 7623 14116
rect 7639 14172 7703 14176
rect 7639 14116 7643 14172
rect 7643 14116 7699 14172
rect 7699 14116 7703 14172
rect 7639 14112 7703 14116
rect 7719 14172 7783 14176
rect 7719 14116 7723 14172
rect 7723 14116 7779 14172
rect 7779 14116 7783 14172
rect 7719 14112 7783 14116
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5847 13628 5911 13632
rect 5847 13572 5851 13628
rect 5851 13572 5907 13628
rect 5907 13572 5911 13628
rect 5847 13568 5911 13572
rect 5927 13628 5991 13632
rect 5927 13572 5931 13628
rect 5931 13572 5987 13628
rect 5987 13572 5991 13628
rect 5927 13568 5991 13572
rect 6007 13628 6071 13632
rect 6007 13572 6011 13628
rect 6011 13572 6067 13628
rect 6067 13572 6071 13628
rect 6007 13568 6071 13572
rect 6087 13628 6151 13632
rect 6087 13572 6091 13628
rect 6091 13572 6147 13628
rect 6147 13572 6151 13628
rect 6087 13568 6151 13572
rect 9111 13628 9175 13632
rect 9111 13572 9115 13628
rect 9115 13572 9171 13628
rect 9171 13572 9175 13628
rect 9111 13568 9175 13572
rect 9191 13628 9255 13632
rect 9191 13572 9195 13628
rect 9195 13572 9251 13628
rect 9251 13572 9255 13628
rect 9191 13568 9255 13572
rect 9271 13628 9335 13632
rect 9271 13572 9275 13628
rect 9275 13572 9331 13628
rect 9331 13572 9335 13628
rect 9271 13568 9335 13572
rect 9351 13628 9415 13632
rect 9351 13572 9355 13628
rect 9355 13572 9411 13628
rect 9411 13572 9415 13628
rect 9351 13568 9415 13572
rect 4215 13084 4279 13088
rect 4215 13028 4219 13084
rect 4219 13028 4275 13084
rect 4275 13028 4279 13084
rect 4215 13024 4279 13028
rect 4295 13084 4359 13088
rect 4295 13028 4299 13084
rect 4299 13028 4355 13084
rect 4355 13028 4359 13084
rect 4295 13024 4359 13028
rect 4375 13084 4439 13088
rect 4375 13028 4379 13084
rect 4379 13028 4435 13084
rect 4435 13028 4439 13084
rect 4375 13024 4439 13028
rect 4455 13084 4519 13088
rect 4455 13028 4459 13084
rect 4459 13028 4515 13084
rect 4515 13028 4519 13084
rect 4455 13024 4519 13028
rect 7479 13084 7543 13088
rect 7479 13028 7483 13084
rect 7483 13028 7539 13084
rect 7539 13028 7543 13084
rect 7479 13024 7543 13028
rect 7559 13084 7623 13088
rect 7559 13028 7563 13084
rect 7563 13028 7619 13084
rect 7619 13028 7623 13084
rect 7559 13024 7623 13028
rect 7639 13084 7703 13088
rect 7639 13028 7643 13084
rect 7643 13028 7699 13084
rect 7699 13028 7703 13084
rect 7639 13024 7703 13028
rect 7719 13084 7783 13088
rect 7719 13028 7723 13084
rect 7723 13028 7779 13084
rect 7779 13028 7783 13084
rect 7719 13024 7783 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5847 12540 5911 12544
rect 5847 12484 5851 12540
rect 5851 12484 5907 12540
rect 5907 12484 5911 12540
rect 5847 12480 5911 12484
rect 5927 12540 5991 12544
rect 5927 12484 5931 12540
rect 5931 12484 5987 12540
rect 5987 12484 5991 12540
rect 5927 12480 5991 12484
rect 6007 12540 6071 12544
rect 6007 12484 6011 12540
rect 6011 12484 6067 12540
rect 6067 12484 6071 12540
rect 6007 12480 6071 12484
rect 6087 12540 6151 12544
rect 6087 12484 6091 12540
rect 6091 12484 6147 12540
rect 6147 12484 6151 12540
rect 6087 12480 6151 12484
rect 9111 12540 9175 12544
rect 9111 12484 9115 12540
rect 9115 12484 9171 12540
rect 9171 12484 9175 12540
rect 9111 12480 9175 12484
rect 9191 12540 9255 12544
rect 9191 12484 9195 12540
rect 9195 12484 9251 12540
rect 9251 12484 9255 12540
rect 9191 12480 9255 12484
rect 9271 12540 9335 12544
rect 9271 12484 9275 12540
rect 9275 12484 9331 12540
rect 9331 12484 9335 12540
rect 9271 12480 9335 12484
rect 9351 12540 9415 12544
rect 9351 12484 9355 12540
rect 9355 12484 9411 12540
rect 9411 12484 9415 12540
rect 9351 12480 9415 12484
rect 4215 11996 4279 12000
rect 4215 11940 4219 11996
rect 4219 11940 4275 11996
rect 4275 11940 4279 11996
rect 4215 11936 4279 11940
rect 4295 11996 4359 12000
rect 4295 11940 4299 11996
rect 4299 11940 4355 11996
rect 4355 11940 4359 11996
rect 4295 11936 4359 11940
rect 4375 11996 4439 12000
rect 4375 11940 4379 11996
rect 4379 11940 4435 11996
rect 4435 11940 4439 11996
rect 4375 11936 4439 11940
rect 4455 11996 4519 12000
rect 4455 11940 4459 11996
rect 4459 11940 4515 11996
rect 4515 11940 4519 11996
rect 4455 11936 4519 11940
rect 7479 11996 7543 12000
rect 7479 11940 7483 11996
rect 7483 11940 7539 11996
rect 7539 11940 7543 11996
rect 7479 11936 7543 11940
rect 7559 11996 7623 12000
rect 7559 11940 7563 11996
rect 7563 11940 7619 11996
rect 7619 11940 7623 11996
rect 7559 11936 7623 11940
rect 7639 11996 7703 12000
rect 7639 11940 7643 11996
rect 7643 11940 7699 11996
rect 7699 11940 7703 11996
rect 7639 11936 7703 11940
rect 7719 11996 7783 12000
rect 7719 11940 7723 11996
rect 7723 11940 7779 11996
rect 7779 11940 7783 11996
rect 7719 11936 7783 11940
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5847 11452 5911 11456
rect 5847 11396 5851 11452
rect 5851 11396 5907 11452
rect 5907 11396 5911 11452
rect 5847 11392 5911 11396
rect 5927 11452 5991 11456
rect 5927 11396 5931 11452
rect 5931 11396 5987 11452
rect 5987 11396 5991 11452
rect 5927 11392 5991 11396
rect 6007 11452 6071 11456
rect 6007 11396 6011 11452
rect 6011 11396 6067 11452
rect 6067 11396 6071 11452
rect 6007 11392 6071 11396
rect 6087 11452 6151 11456
rect 6087 11396 6091 11452
rect 6091 11396 6147 11452
rect 6147 11396 6151 11452
rect 6087 11392 6151 11396
rect 9111 11452 9175 11456
rect 9111 11396 9115 11452
rect 9115 11396 9171 11452
rect 9171 11396 9175 11452
rect 9111 11392 9175 11396
rect 9191 11452 9255 11456
rect 9191 11396 9195 11452
rect 9195 11396 9251 11452
rect 9251 11396 9255 11452
rect 9191 11392 9255 11396
rect 9271 11452 9335 11456
rect 9271 11396 9275 11452
rect 9275 11396 9331 11452
rect 9331 11396 9335 11452
rect 9271 11392 9335 11396
rect 9351 11452 9415 11456
rect 9351 11396 9355 11452
rect 9355 11396 9411 11452
rect 9411 11396 9415 11452
rect 9351 11392 9415 11396
rect 4215 10908 4279 10912
rect 4215 10852 4219 10908
rect 4219 10852 4275 10908
rect 4275 10852 4279 10908
rect 4215 10848 4279 10852
rect 4295 10908 4359 10912
rect 4295 10852 4299 10908
rect 4299 10852 4355 10908
rect 4355 10852 4359 10908
rect 4295 10848 4359 10852
rect 4375 10908 4439 10912
rect 4375 10852 4379 10908
rect 4379 10852 4435 10908
rect 4435 10852 4439 10908
rect 4375 10848 4439 10852
rect 4455 10908 4519 10912
rect 4455 10852 4459 10908
rect 4459 10852 4515 10908
rect 4515 10852 4519 10908
rect 4455 10848 4519 10852
rect 7479 10908 7543 10912
rect 7479 10852 7483 10908
rect 7483 10852 7539 10908
rect 7539 10852 7543 10908
rect 7479 10848 7543 10852
rect 7559 10908 7623 10912
rect 7559 10852 7563 10908
rect 7563 10852 7619 10908
rect 7619 10852 7623 10908
rect 7559 10848 7623 10852
rect 7639 10908 7703 10912
rect 7639 10852 7643 10908
rect 7643 10852 7699 10908
rect 7699 10852 7703 10908
rect 7639 10848 7703 10852
rect 7719 10908 7783 10912
rect 7719 10852 7723 10908
rect 7723 10852 7779 10908
rect 7779 10852 7783 10908
rect 7719 10848 7783 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5847 10364 5911 10368
rect 5847 10308 5851 10364
rect 5851 10308 5907 10364
rect 5907 10308 5911 10364
rect 5847 10304 5911 10308
rect 5927 10364 5991 10368
rect 5927 10308 5931 10364
rect 5931 10308 5987 10364
rect 5987 10308 5991 10364
rect 5927 10304 5991 10308
rect 6007 10364 6071 10368
rect 6007 10308 6011 10364
rect 6011 10308 6067 10364
rect 6067 10308 6071 10364
rect 6007 10304 6071 10308
rect 6087 10364 6151 10368
rect 6087 10308 6091 10364
rect 6091 10308 6147 10364
rect 6147 10308 6151 10364
rect 6087 10304 6151 10308
rect 9111 10364 9175 10368
rect 9111 10308 9115 10364
rect 9115 10308 9171 10364
rect 9171 10308 9175 10364
rect 9111 10304 9175 10308
rect 9191 10364 9255 10368
rect 9191 10308 9195 10364
rect 9195 10308 9251 10364
rect 9251 10308 9255 10364
rect 9191 10304 9255 10308
rect 9271 10364 9335 10368
rect 9271 10308 9275 10364
rect 9275 10308 9331 10364
rect 9331 10308 9335 10364
rect 9271 10304 9335 10308
rect 9351 10364 9415 10368
rect 9351 10308 9355 10364
rect 9355 10308 9411 10364
rect 9411 10308 9415 10364
rect 9351 10304 9415 10308
rect 4215 9820 4279 9824
rect 4215 9764 4219 9820
rect 4219 9764 4275 9820
rect 4275 9764 4279 9820
rect 4215 9760 4279 9764
rect 4295 9820 4359 9824
rect 4295 9764 4299 9820
rect 4299 9764 4355 9820
rect 4355 9764 4359 9820
rect 4295 9760 4359 9764
rect 4375 9820 4439 9824
rect 4375 9764 4379 9820
rect 4379 9764 4435 9820
rect 4435 9764 4439 9820
rect 4375 9760 4439 9764
rect 4455 9820 4519 9824
rect 4455 9764 4459 9820
rect 4459 9764 4515 9820
rect 4515 9764 4519 9820
rect 4455 9760 4519 9764
rect 7479 9820 7543 9824
rect 7479 9764 7483 9820
rect 7483 9764 7539 9820
rect 7539 9764 7543 9820
rect 7479 9760 7543 9764
rect 7559 9820 7623 9824
rect 7559 9764 7563 9820
rect 7563 9764 7619 9820
rect 7619 9764 7623 9820
rect 7559 9760 7623 9764
rect 7639 9820 7703 9824
rect 7639 9764 7643 9820
rect 7643 9764 7699 9820
rect 7699 9764 7703 9820
rect 7639 9760 7703 9764
rect 7719 9820 7783 9824
rect 7719 9764 7723 9820
rect 7723 9764 7779 9820
rect 7779 9764 7783 9820
rect 7719 9760 7783 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5847 9276 5911 9280
rect 5847 9220 5851 9276
rect 5851 9220 5907 9276
rect 5907 9220 5911 9276
rect 5847 9216 5911 9220
rect 5927 9276 5991 9280
rect 5927 9220 5931 9276
rect 5931 9220 5987 9276
rect 5987 9220 5991 9276
rect 5927 9216 5991 9220
rect 6007 9276 6071 9280
rect 6007 9220 6011 9276
rect 6011 9220 6067 9276
rect 6067 9220 6071 9276
rect 6007 9216 6071 9220
rect 6087 9276 6151 9280
rect 6087 9220 6091 9276
rect 6091 9220 6147 9276
rect 6147 9220 6151 9276
rect 6087 9216 6151 9220
rect 9111 9276 9175 9280
rect 9111 9220 9115 9276
rect 9115 9220 9171 9276
rect 9171 9220 9175 9276
rect 9111 9216 9175 9220
rect 9191 9276 9255 9280
rect 9191 9220 9195 9276
rect 9195 9220 9251 9276
rect 9251 9220 9255 9276
rect 9191 9216 9255 9220
rect 9271 9276 9335 9280
rect 9271 9220 9275 9276
rect 9275 9220 9331 9276
rect 9331 9220 9335 9276
rect 9271 9216 9335 9220
rect 9351 9276 9415 9280
rect 9351 9220 9355 9276
rect 9355 9220 9411 9276
rect 9411 9220 9415 9276
rect 9351 9216 9415 9220
rect 4215 8732 4279 8736
rect 4215 8676 4219 8732
rect 4219 8676 4275 8732
rect 4275 8676 4279 8732
rect 4215 8672 4279 8676
rect 4295 8732 4359 8736
rect 4295 8676 4299 8732
rect 4299 8676 4355 8732
rect 4355 8676 4359 8732
rect 4295 8672 4359 8676
rect 4375 8732 4439 8736
rect 4375 8676 4379 8732
rect 4379 8676 4435 8732
rect 4435 8676 4439 8732
rect 4375 8672 4439 8676
rect 4455 8732 4519 8736
rect 4455 8676 4459 8732
rect 4459 8676 4515 8732
rect 4515 8676 4519 8732
rect 4455 8672 4519 8676
rect 7479 8732 7543 8736
rect 7479 8676 7483 8732
rect 7483 8676 7539 8732
rect 7539 8676 7543 8732
rect 7479 8672 7543 8676
rect 7559 8732 7623 8736
rect 7559 8676 7563 8732
rect 7563 8676 7619 8732
rect 7619 8676 7623 8732
rect 7559 8672 7623 8676
rect 7639 8732 7703 8736
rect 7639 8676 7643 8732
rect 7643 8676 7699 8732
rect 7699 8676 7703 8732
rect 7639 8672 7703 8676
rect 7719 8732 7783 8736
rect 7719 8676 7723 8732
rect 7723 8676 7779 8732
rect 7779 8676 7783 8732
rect 7719 8672 7783 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5847 8188 5911 8192
rect 5847 8132 5851 8188
rect 5851 8132 5907 8188
rect 5907 8132 5911 8188
rect 5847 8128 5911 8132
rect 5927 8188 5991 8192
rect 5927 8132 5931 8188
rect 5931 8132 5987 8188
rect 5987 8132 5991 8188
rect 5927 8128 5991 8132
rect 6007 8188 6071 8192
rect 6007 8132 6011 8188
rect 6011 8132 6067 8188
rect 6067 8132 6071 8188
rect 6007 8128 6071 8132
rect 6087 8188 6151 8192
rect 6087 8132 6091 8188
rect 6091 8132 6147 8188
rect 6147 8132 6151 8188
rect 6087 8128 6151 8132
rect 9111 8188 9175 8192
rect 9111 8132 9115 8188
rect 9115 8132 9171 8188
rect 9171 8132 9175 8188
rect 9111 8128 9175 8132
rect 9191 8188 9255 8192
rect 9191 8132 9195 8188
rect 9195 8132 9251 8188
rect 9251 8132 9255 8188
rect 9191 8128 9255 8132
rect 9271 8188 9335 8192
rect 9271 8132 9275 8188
rect 9275 8132 9331 8188
rect 9331 8132 9335 8188
rect 9271 8128 9335 8132
rect 9351 8188 9415 8192
rect 9351 8132 9355 8188
rect 9355 8132 9411 8188
rect 9411 8132 9415 8188
rect 9351 8128 9415 8132
rect 4215 7644 4279 7648
rect 4215 7588 4219 7644
rect 4219 7588 4275 7644
rect 4275 7588 4279 7644
rect 4215 7584 4279 7588
rect 4295 7644 4359 7648
rect 4295 7588 4299 7644
rect 4299 7588 4355 7644
rect 4355 7588 4359 7644
rect 4295 7584 4359 7588
rect 4375 7644 4439 7648
rect 4375 7588 4379 7644
rect 4379 7588 4435 7644
rect 4435 7588 4439 7644
rect 4375 7584 4439 7588
rect 4455 7644 4519 7648
rect 4455 7588 4459 7644
rect 4459 7588 4515 7644
rect 4515 7588 4519 7644
rect 4455 7584 4519 7588
rect 7479 7644 7543 7648
rect 7479 7588 7483 7644
rect 7483 7588 7539 7644
rect 7539 7588 7543 7644
rect 7479 7584 7543 7588
rect 7559 7644 7623 7648
rect 7559 7588 7563 7644
rect 7563 7588 7619 7644
rect 7619 7588 7623 7644
rect 7559 7584 7623 7588
rect 7639 7644 7703 7648
rect 7639 7588 7643 7644
rect 7643 7588 7699 7644
rect 7699 7588 7703 7644
rect 7639 7584 7703 7588
rect 7719 7644 7783 7648
rect 7719 7588 7723 7644
rect 7723 7588 7779 7644
rect 7779 7588 7783 7644
rect 7719 7584 7783 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5847 7100 5911 7104
rect 5847 7044 5851 7100
rect 5851 7044 5907 7100
rect 5907 7044 5911 7100
rect 5847 7040 5911 7044
rect 5927 7100 5991 7104
rect 5927 7044 5931 7100
rect 5931 7044 5987 7100
rect 5987 7044 5991 7100
rect 5927 7040 5991 7044
rect 6007 7100 6071 7104
rect 6007 7044 6011 7100
rect 6011 7044 6067 7100
rect 6067 7044 6071 7100
rect 6007 7040 6071 7044
rect 6087 7100 6151 7104
rect 6087 7044 6091 7100
rect 6091 7044 6147 7100
rect 6147 7044 6151 7100
rect 6087 7040 6151 7044
rect 9111 7100 9175 7104
rect 9111 7044 9115 7100
rect 9115 7044 9171 7100
rect 9171 7044 9175 7100
rect 9111 7040 9175 7044
rect 9191 7100 9255 7104
rect 9191 7044 9195 7100
rect 9195 7044 9251 7100
rect 9251 7044 9255 7100
rect 9191 7040 9255 7044
rect 9271 7100 9335 7104
rect 9271 7044 9275 7100
rect 9275 7044 9331 7100
rect 9331 7044 9335 7100
rect 9271 7040 9335 7044
rect 9351 7100 9415 7104
rect 9351 7044 9355 7100
rect 9355 7044 9411 7100
rect 9411 7044 9415 7100
rect 9351 7040 9415 7044
rect 4215 6556 4279 6560
rect 4215 6500 4219 6556
rect 4219 6500 4275 6556
rect 4275 6500 4279 6556
rect 4215 6496 4279 6500
rect 4295 6556 4359 6560
rect 4295 6500 4299 6556
rect 4299 6500 4355 6556
rect 4355 6500 4359 6556
rect 4295 6496 4359 6500
rect 4375 6556 4439 6560
rect 4375 6500 4379 6556
rect 4379 6500 4435 6556
rect 4435 6500 4439 6556
rect 4375 6496 4439 6500
rect 4455 6556 4519 6560
rect 4455 6500 4459 6556
rect 4459 6500 4515 6556
rect 4515 6500 4519 6556
rect 4455 6496 4519 6500
rect 7479 6556 7543 6560
rect 7479 6500 7483 6556
rect 7483 6500 7539 6556
rect 7539 6500 7543 6556
rect 7479 6496 7543 6500
rect 7559 6556 7623 6560
rect 7559 6500 7563 6556
rect 7563 6500 7619 6556
rect 7619 6500 7623 6556
rect 7559 6496 7623 6500
rect 7639 6556 7703 6560
rect 7639 6500 7643 6556
rect 7643 6500 7699 6556
rect 7699 6500 7703 6556
rect 7639 6496 7703 6500
rect 7719 6556 7783 6560
rect 7719 6500 7723 6556
rect 7723 6500 7779 6556
rect 7779 6500 7783 6556
rect 7719 6496 7783 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5847 6012 5911 6016
rect 5847 5956 5851 6012
rect 5851 5956 5907 6012
rect 5907 5956 5911 6012
rect 5847 5952 5911 5956
rect 5927 6012 5991 6016
rect 5927 5956 5931 6012
rect 5931 5956 5987 6012
rect 5987 5956 5991 6012
rect 5927 5952 5991 5956
rect 6007 6012 6071 6016
rect 6007 5956 6011 6012
rect 6011 5956 6067 6012
rect 6067 5956 6071 6012
rect 6007 5952 6071 5956
rect 6087 6012 6151 6016
rect 6087 5956 6091 6012
rect 6091 5956 6147 6012
rect 6147 5956 6151 6012
rect 6087 5952 6151 5956
rect 9111 6012 9175 6016
rect 9111 5956 9115 6012
rect 9115 5956 9171 6012
rect 9171 5956 9175 6012
rect 9111 5952 9175 5956
rect 9191 6012 9255 6016
rect 9191 5956 9195 6012
rect 9195 5956 9251 6012
rect 9251 5956 9255 6012
rect 9191 5952 9255 5956
rect 9271 6012 9335 6016
rect 9271 5956 9275 6012
rect 9275 5956 9331 6012
rect 9331 5956 9335 6012
rect 9271 5952 9335 5956
rect 9351 6012 9415 6016
rect 9351 5956 9355 6012
rect 9355 5956 9411 6012
rect 9411 5956 9415 6012
rect 9351 5952 9415 5956
rect 4215 5468 4279 5472
rect 4215 5412 4219 5468
rect 4219 5412 4275 5468
rect 4275 5412 4279 5468
rect 4215 5408 4279 5412
rect 4295 5468 4359 5472
rect 4295 5412 4299 5468
rect 4299 5412 4355 5468
rect 4355 5412 4359 5468
rect 4295 5408 4359 5412
rect 4375 5468 4439 5472
rect 4375 5412 4379 5468
rect 4379 5412 4435 5468
rect 4435 5412 4439 5468
rect 4375 5408 4439 5412
rect 4455 5468 4519 5472
rect 4455 5412 4459 5468
rect 4459 5412 4515 5468
rect 4515 5412 4519 5468
rect 4455 5408 4519 5412
rect 7479 5468 7543 5472
rect 7479 5412 7483 5468
rect 7483 5412 7539 5468
rect 7539 5412 7543 5468
rect 7479 5408 7543 5412
rect 7559 5468 7623 5472
rect 7559 5412 7563 5468
rect 7563 5412 7619 5468
rect 7619 5412 7623 5468
rect 7559 5408 7623 5412
rect 7639 5468 7703 5472
rect 7639 5412 7643 5468
rect 7643 5412 7699 5468
rect 7699 5412 7703 5468
rect 7639 5408 7703 5412
rect 7719 5468 7783 5472
rect 7719 5412 7723 5468
rect 7723 5412 7779 5468
rect 7779 5412 7783 5468
rect 7719 5408 7783 5412
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5847 4924 5911 4928
rect 5847 4868 5851 4924
rect 5851 4868 5907 4924
rect 5907 4868 5911 4924
rect 5847 4864 5911 4868
rect 5927 4924 5991 4928
rect 5927 4868 5931 4924
rect 5931 4868 5987 4924
rect 5987 4868 5991 4924
rect 5927 4864 5991 4868
rect 6007 4924 6071 4928
rect 6007 4868 6011 4924
rect 6011 4868 6067 4924
rect 6067 4868 6071 4924
rect 6007 4864 6071 4868
rect 6087 4924 6151 4928
rect 6087 4868 6091 4924
rect 6091 4868 6147 4924
rect 6147 4868 6151 4924
rect 6087 4864 6151 4868
rect 9111 4924 9175 4928
rect 9111 4868 9115 4924
rect 9115 4868 9171 4924
rect 9171 4868 9175 4924
rect 9111 4864 9175 4868
rect 9191 4924 9255 4928
rect 9191 4868 9195 4924
rect 9195 4868 9251 4924
rect 9251 4868 9255 4924
rect 9191 4864 9255 4868
rect 9271 4924 9335 4928
rect 9271 4868 9275 4924
rect 9275 4868 9331 4924
rect 9331 4868 9335 4924
rect 9271 4864 9335 4868
rect 9351 4924 9415 4928
rect 9351 4868 9355 4924
rect 9355 4868 9411 4924
rect 9411 4868 9415 4924
rect 9351 4864 9415 4868
rect 4215 4380 4279 4384
rect 4215 4324 4219 4380
rect 4219 4324 4275 4380
rect 4275 4324 4279 4380
rect 4215 4320 4279 4324
rect 4295 4380 4359 4384
rect 4295 4324 4299 4380
rect 4299 4324 4355 4380
rect 4355 4324 4359 4380
rect 4295 4320 4359 4324
rect 4375 4380 4439 4384
rect 4375 4324 4379 4380
rect 4379 4324 4435 4380
rect 4435 4324 4439 4380
rect 4375 4320 4439 4324
rect 4455 4380 4519 4384
rect 4455 4324 4459 4380
rect 4459 4324 4515 4380
rect 4515 4324 4519 4380
rect 4455 4320 4519 4324
rect 7479 4380 7543 4384
rect 7479 4324 7483 4380
rect 7483 4324 7539 4380
rect 7539 4324 7543 4380
rect 7479 4320 7543 4324
rect 7559 4380 7623 4384
rect 7559 4324 7563 4380
rect 7563 4324 7619 4380
rect 7619 4324 7623 4380
rect 7559 4320 7623 4324
rect 7639 4380 7703 4384
rect 7639 4324 7643 4380
rect 7643 4324 7699 4380
rect 7699 4324 7703 4380
rect 7639 4320 7703 4324
rect 7719 4380 7783 4384
rect 7719 4324 7723 4380
rect 7723 4324 7779 4380
rect 7779 4324 7783 4380
rect 7719 4320 7783 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5847 3836 5911 3840
rect 5847 3780 5851 3836
rect 5851 3780 5907 3836
rect 5907 3780 5911 3836
rect 5847 3776 5911 3780
rect 5927 3836 5991 3840
rect 5927 3780 5931 3836
rect 5931 3780 5987 3836
rect 5987 3780 5991 3836
rect 5927 3776 5991 3780
rect 6007 3836 6071 3840
rect 6007 3780 6011 3836
rect 6011 3780 6067 3836
rect 6067 3780 6071 3836
rect 6007 3776 6071 3780
rect 6087 3836 6151 3840
rect 6087 3780 6091 3836
rect 6091 3780 6147 3836
rect 6147 3780 6151 3836
rect 6087 3776 6151 3780
rect 9111 3836 9175 3840
rect 9111 3780 9115 3836
rect 9115 3780 9171 3836
rect 9171 3780 9175 3836
rect 9111 3776 9175 3780
rect 9191 3836 9255 3840
rect 9191 3780 9195 3836
rect 9195 3780 9251 3836
rect 9251 3780 9255 3836
rect 9191 3776 9255 3780
rect 9271 3836 9335 3840
rect 9271 3780 9275 3836
rect 9275 3780 9331 3836
rect 9331 3780 9335 3836
rect 9271 3776 9335 3780
rect 9351 3836 9415 3840
rect 9351 3780 9355 3836
rect 9355 3780 9411 3836
rect 9411 3780 9415 3836
rect 9351 3776 9415 3780
rect 4215 3292 4279 3296
rect 4215 3236 4219 3292
rect 4219 3236 4275 3292
rect 4275 3236 4279 3292
rect 4215 3232 4279 3236
rect 4295 3292 4359 3296
rect 4295 3236 4299 3292
rect 4299 3236 4355 3292
rect 4355 3236 4359 3292
rect 4295 3232 4359 3236
rect 4375 3292 4439 3296
rect 4375 3236 4379 3292
rect 4379 3236 4435 3292
rect 4435 3236 4439 3292
rect 4375 3232 4439 3236
rect 4455 3292 4519 3296
rect 4455 3236 4459 3292
rect 4459 3236 4515 3292
rect 4515 3236 4519 3292
rect 4455 3232 4519 3236
rect 7479 3292 7543 3296
rect 7479 3236 7483 3292
rect 7483 3236 7539 3292
rect 7539 3236 7543 3292
rect 7479 3232 7543 3236
rect 7559 3292 7623 3296
rect 7559 3236 7563 3292
rect 7563 3236 7619 3292
rect 7619 3236 7623 3292
rect 7559 3232 7623 3236
rect 7639 3292 7703 3296
rect 7639 3236 7643 3292
rect 7643 3236 7699 3292
rect 7699 3236 7703 3292
rect 7639 3232 7703 3236
rect 7719 3292 7783 3296
rect 7719 3236 7723 3292
rect 7723 3236 7779 3292
rect 7779 3236 7783 3292
rect 7719 3232 7783 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5847 2748 5911 2752
rect 5847 2692 5851 2748
rect 5851 2692 5907 2748
rect 5907 2692 5911 2748
rect 5847 2688 5911 2692
rect 5927 2748 5991 2752
rect 5927 2692 5931 2748
rect 5931 2692 5987 2748
rect 5987 2692 5991 2748
rect 5927 2688 5991 2692
rect 6007 2748 6071 2752
rect 6007 2692 6011 2748
rect 6011 2692 6067 2748
rect 6067 2692 6071 2748
rect 6007 2688 6071 2692
rect 6087 2748 6151 2752
rect 6087 2692 6091 2748
rect 6091 2692 6147 2748
rect 6147 2692 6151 2748
rect 6087 2688 6151 2692
rect 9111 2748 9175 2752
rect 9111 2692 9115 2748
rect 9115 2692 9171 2748
rect 9171 2692 9175 2748
rect 9111 2688 9175 2692
rect 9191 2748 9255 2752
rect 9191 2692 9195 2748
rect 9195 2692 9251 2748
rect 9251 2692 9255 2748
rect 9191 2688 9255 2692
rect 9271 2748 9335 2752
rect 9271 2692 9275 2748
rect 9275 2692 9331 2748
rect 9331 2692 9335 2748
rect 9271 2688 9335 2692
rect 9351 2748 9415 2752
rect 9351 2692 9355 2748
rect 9355 2692 9411 2748
rect 9411 2692 9415 2748
rect 9351 2688 9415 2692
rect 4215 2204 4279 2208
rect 4215 2148 4219 2204
rect 4219 2148 4275 2204
rect 4275 2148 4279 2204
rect 4215 2144 4279 2148
rect 4295 2204 4359 2208
rect 4295 2148 4299 2204
rect 4299 2148 4355 2204
rect 4355 2148 4359 2204
rect 4295 2144 4359 2148
rect 4375 2204 4439 2208
rect 4375 2148 4379 2204
rect 4379 2148 4435 2204
rect 4435 2148 4439 2204
rect 4375 2144 4439 2148
rect 4455 2204 4519 2208
rect 4455 2148 4459 2204
rect 4459 2148 4515 2204
rect 4515 2148 4519 2204
rect 4455 2144 4519 2148
rect 7479 2204 7543 2208
rect 7479 2148 7483 2204
rect 7483 2148 7539 2204
rect 7539 2148 7543 2204
rect 7479 2144 7543 2148
rect 7559 2204 7623 2208
rect 7559 2148 7563 2204
rect 7563 2148 7619 2204
rect 7619 2148 7623 2204
rect 7559 2144 7623 2148
rect 7639 2204 7703 2208
rect 7639 2148 7643 2204
rect 7643 2148 7699 2204
rect 7699 2148 7703 2204
rect 7639 2144 7703 2148
rect 7719 2204 7783 2208
rect 7719 2148 7723 2204
rect 7723 2148 7779 2204
rect 7779 2148 7783 2204
rect 7719 2144 7783 2148
<< metal4 >>
rect 2575 77824 2896 77840
rect 2575 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2575 76736 2896 77760
rect 2575 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2575 75648 2896 76672
rect 2575 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2575 74560 2896 75584
rect 2575 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2575 73472 2896 74496
rect 2575 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2575 72384 2896 73408
rect 2575 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2575 71296 2896 72320
rect 2575 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2575 70208 2896 71232
rect 2575 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2575 69120 2896 70144
rect 2575 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2575 68032 2896 69056
rect 2575 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2575 66944 2896 67968
rect 2575 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2083 66468 2149 66469
rect 2083 66404 2084 66468
rect 2148 66404 2149 66468
rect 2083 66403 2149 66404
rect 1899 64972 1965 64973
rect 1899 64908 1900 64972
rect 1964 64908 1965 64972
rect 1899 64907 1965 64908
rect 1715 59668 1781 59669
rect 1715 59604 1716 59668
rect 1780 59604 1781 59668
rect 1715 59603 1781 59604
rect 1718 51917 1778 59603
rect 1902 58853 1962 64907
rect 2086 60757 2146 66403
rect 2575 65856 2896 66880
rect 2575 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2575 64768 2896 65792
rect 2575 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2575 63680 2896 64704
rect 2575 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2575 62592 2896 63616
rect 2575 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2575 61504 2896 62528
rect 2575 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2267 60892 2333 60893
rect 2267 60828 2268 60892
rect 2332 60828 2333 60892
rect 2267 60827 2333 60828
rect 2083 60756 2149 60757
rect 2083 60692 2084 60756
rect 2148 60692 2149 60756
rect 2083 60691 2149 60692
rect 2270 60213 2330 60827
rect 2575 60416 2896 61440
rect 2575 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2267 60212 2333 60213
rect 2267 60148 2268 60212
rect 2332 60148 2333 60212
rect 2267 60147 2333 60148
rect 2575 59328 2896 60352
rect 2575 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 1899 58852 1965 58853
rect 1899 58788 1900 58852
rect 1964 58788 1965 58852
rect 1899 58787 1965 58788
rect 2575 58240 2896 59264
rect 2575 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2575 57152 2896 58176
rect 4207 77280 4527 77840
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 76192 4527 77216
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 75104 4527 76128
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 74016 4527 75040
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 72928 4527 73952
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 71840 4527 72864
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 70752 4527 71776
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 69664 4527 70688
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 68576 4527 69600
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 67488 4527 68512
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 66400 4527 67424
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 65312 4527 66336
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 64224 4527 65248
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 63136 4527 64160
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 62048 4527 63072
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 60960 4527 61984
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 59872 4527 60896
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 58784 4527 59808
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 3187 57900 3253 57901
rect 3187 57836 3188 57900
rect 3252 57836 3253 57900
rect 3187 57835 3253 57836
rect 2575 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2575 56064 2896 57088
rect 2575 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2575 54976 2896 56000
rect 2575 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2575 53888 2896 54912
rect 2575 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2575 52800 2896 53824
rect 2575 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 1715 51916 1781 51917
rect 1715 51852 1716 51916
rect 1780 51852 1781 51916
rect 1715 51851 1781 51852
rect 2575 51712 2896 52736
rect 2575 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2575 50624 2896 51648
rect 2575 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2575 49536 2896 50560
rect 3190 50421 3250 57835
rect 4207 57696 4527 58720
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 3371 56948 3437 56949
rect 3371 56884 3372 56948
rect 3436 56884 3437 56948
rect 3371 56883 3437 56884
rect 3187 50420 3253 50421
rect 3187 50356 3188 50420
rect 3252 50356 3253 50420
rect 3187 50355 3253 50356
rect 2575 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2575 48448 2896 49472
rect 2575 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 1899 48380 1965 48381
rect 1899 48316 1900 48380
rect 1964 48316 1965 48380
rect 1899 48315 1965 48316
rect 1902 40085 1962 48315
rect 2575 47360 2896 48384
rect 3374 48381 3434 56883
rect 4207 56608 4527 57632
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 55520 4527 56544
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 54432 4527 55456
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 53344 4527 54368
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 52256 4527 53280
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 51168 4527 52192
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 50080 4527 51104
rect 5839 77824 6159 77840
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 76736 6159 77760
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 75648 6159 76672
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 74560 6159 75584
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 73472 6159 74496
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 72384 6159 73408
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 71296 6159 72320
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 70208 6159 71232
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 69120 6159 70144
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 68032 6159 69056
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 66944 6159 67968
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 65856 6159 66880
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 64768 6159 65792
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 63680 6159 64704
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 62592 6159 63616
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 61504 6159 62528
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 60416 6159 61440
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 59328 6159 60352
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 58240 6159 59264
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 57152 6159 58176
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 56064 6159 57088
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 54976 6159 56000
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 53888 6159 54912
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 52800 6159 53824
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 51712 6159 52736
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 50624 6159 51648
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 4659 50420 4725 50421
rect 4659 50356 4660 50420
rect 4724 50356 4725 50420
rect 4659 50355 4725 50356
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 48992 4527 50016
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 3371 48380 3437 48381
rect 3371 48316 3372 48380
rect 3436 48316 3437 48380
rect 3371 48315 3437 48316
rect 4207 47904 4527 48928
rect 4662 48789 4722 50355
rect 5839 49536 6159 50560
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 4659 48788 4725 48789
rect 4659 48724 4660 48788
rect 4724 48724 4725 48788
rect 4659 48723 4725 48724
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 3003 47836 3069 47837
rect 3003 47772 3004 47836
rect 3068 47772 3069 47836
rect 3003 47771 3069 47772
rect 2575 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2083 47156 2149 47157
rect 2083 47092 2084 47156
rect 2148 47092 2149 47156
rect 2083 47091 2149 47092
rect 2086 40901 2146 47091
rect 2575 46272 2896 47296
rect 3006 46477 3066 47771
rect 4207 46816 4527 47840
rect 5839 48448 6159 49472
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 4659 47564 4725 47565
rect 4659 47500 4660 47564
rect 4724 47500 4725 47564
rect 4659 47499 4725 47500
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 3003 46476 3069 46477
rect 3003 46412 3004 46476
rect 3068 46412 3069 46476
rect 3003 46411 3069 46412
rect 2575 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2575 45184 2896 46208
rect 2575 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2575 44096 2896 45120
rect 3006 44437 3066 46411
rect 4207 45728 4527 46752
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 44640 4527 45664
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 3003 44436 3069 44437
rect 3003 44372 3004 44436
rect 3068 44372 3069 44436
rect 3003 44371 3069 44372
rect 2575 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2575 43008 2896 44032
rect 2575 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2575 41920 2896 42944
rect 2575 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2267 41172 2333 41173
rect 2267 41108 2268 41172
rect 2332 41108 2333 41172
rect 2267 41107 2333 41108
rect 2083 40900 2149 40901
rect 2083 40836 2084 40900
rect 2148 40836 2149 40900
rect 2083 40835 2149 40836
rect 1899 40084 1965 40085
rect 1899 40020 1900 40084
rect 1964 40020 1965 40084
rect 1899 40019 1965 40020
rect 1899 31924 1965 31925
rect 1899 31860 1900 31924
rect 1964 31860 1965 31924
rect 1899 31859 1965 31860
rect 1902 28117 1962 31859
rect 2270 31789 2330 41107
rect 2575 40832 2896 41856
rect 4207 43552 4527 44576
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 42464 4527 43488
rect 4662 42533 4722 47499
rect 5839 47360 6159 48384
rect 7471 77280 7791 77840
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 76192 7791 77216
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 75104 7791 76128
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 74016 7791 75040
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 72928 7791 73952
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 71840 7791 72864
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 70752 7791 71776
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 69664 7791 70688
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 68576 7791 69600
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 67488 7791 68512
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 66400 7791 67424
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 65312 7791 66336
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 64224 7791 65248
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 63136 7791 64160
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 62048 7791 63072
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 60960 7791 61984
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 59872 7791 60896
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 58784 7791 59808
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 57696 7791 58720
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 56608 7791 57632
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 55520 7791 56544
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 54432 7791 55456
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 53344 7791 54368
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 52256 7791 53280
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 51168 7791 52192
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 50080 7791 51104
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 48992 7791 50016
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 47904 7791 48928
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 6315 47564 6381 47565
rect 6315 47500 6316 47564
rect 6380 47500 6381 47564
rect 6315 47499 6381 47500
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 46272 6159 47296
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 45184 6159 46208
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 44096 6159 45120
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 43008 6159 44032
rect 6318 43757 6378 47499
rect 7471 46816 7791 47840
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 45728 7791 46752
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 44640 7791 45664
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 6315 43756 6381 43757
rect 6315 43692 6316 43756
rect 6380 43692 6381 43756
rect 6315 43691 6381 43692
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 4659 42532 4725 42533
rect 4659 42468 4660 42532
rect 4724 42468 4725 42532
rect 4659 42467 4725 42468
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 3003 41580 3069 41581
rect 3003 41516 3004 41580
rect 3068 41516 3069 41580
rect 3003 41515 3069 41516
rect 3006 41173 3066 41515
rect 4207 41376 4527 42400
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 3003 41172 3069 41173
rect 3003 41108 3004 41172
rect 3068 41108 3069 41172
rect 3003 41107 3069 41108
rect 2575 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2575 39744 2896 40768
rect 2575 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2575 38656 2896 39680
rect 2575 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2575 37568 2896 38592
rect 4207 40288 4527 41312
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 39200 4527 40224
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 3739 38316 3805 38317
rect 3739 38252 3740 38316
rect 3804 38252 3805 38316
rect 3739 38251 3805 38252
rect 2575 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2575 36480 2896 37504
rect 3371 37364 3437 37365
rect 3371 37300 3372 37364
rect 3436 37300 3437 37364
rect 3371 37299 3437 37300
rect 2575 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2575 35392 2896 36416
rect 2575 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2575 34304 2896 35328
rect 2575 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2575 33216 2896 34240
rect 3374 33557 3434 37299
rect 3371 33556 3437 33557
rect 3371 33492 3372 33556
rect 3436 33492 3437 33556
rect 3371 33491 3437 33492
rect 2575 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2575 32128 2896 33152
rect 2575 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2267 31788 2333 31789
rect 2267 31724 2268 31788
rect 2332 31724 2333 31788
rect 2267 31723 2333 31724
rect 2575 31040 2896 32064
rect 3003 32060 3069 32061
rect 3003 31996 3004 32060
rect 3068 31996 3069 32060
rect 3003 31995 3069 31996
rect 2575 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2575 29952 2896 30976
rect 2575 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2575 28864 2896 29888
rect 2575 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 1899 28116 1965 28117
rect 1899 28052 1900 28116
rect 1964 28052 1965 28116
rect 1899 28051 1965 28052
rect 2575 27776 2896 28800
rect 2575 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2575 26688 2896 27712
rect 3006 27573 3066 31995
rect 3742 30157 3802 38251
rect 4207 38112 4527 39136
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 37024 4527 38048
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 35936 4527 36960
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 34848 4527 35872
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 33760 4527 34784
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 32672 4527 33696
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 31584 4527 32608
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 30496 4527 31520
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 3739 30156 3805 30157
rect 3739 30092 3740 30156
rect 3804 30092 3805 30156
rect 3739 30091 3805 30092
rect 4207 29408 4527 30432
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 3187 28796 3253 28797
rect 3187 28732 3188 28796
rect 3252 28732 3253 28796
rect 3187 28731 3253 28732
rect 3003 27572 3069 27573
rect 3003 27508 3004 27572
rect 3068 27508 3069 27572
rect 3003 27507 3069 27508
rect 2575 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2575 25600 2896 26624
rect 2575 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2575 24512 2896 25536
rect 2575 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2575 23424 2896 24448
rect 2575 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2575 22336 2896 23360
rect 2575 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2575 21248 2896 22272
rect 3190 21997 3250 28731
rect 4207 28320 4527 29344
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 27232 4527 28256
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 26144 4527 27168
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 25056 4527 26080
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 23968 4527 24992
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 22880 4527 23904
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 3187 21996 3253 21997
rect 3187 21932 3188 21996
rect 3252 21932 3253 21996
rect 3187 21931 3253 21932
rect 2575 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2575 20160 2896 21184
rect 2575 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2575 19072 2896 20096
rect 2575 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2575 17984 2896 19008
rect 2575 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2575 16896 2896 17920
rect 2575 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2575 15808 2896 16832
rect 2575 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2575 14720 2896 15744
rect 2575 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2575 13632 2896 14656
rect 2575 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2575 12544 2896 13568
rect 2575 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2575 11456 2896 12480
rect 2575 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2575 10368 2896 11392
rect 2575 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2575 9280 2896 10304
rect 2575 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2575 8192 2896 9216
rect 2575 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2575 7104 2896 8128
rect 2575 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2575 6016 2896 7040
rect 2575 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2575 4928 2896 5952
rect 2575 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2575 3840 2896 4864
rect 2575 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2575 2752 2896 3776
rect 2575 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2575 2128 2896 2688
rect 4207 21792 4527 22816
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 20704 4527 21728
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 19616 4527 20640
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 18528 4527 19552
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 17440 4527 18464
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 16352 4527 17376
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 15264 4527 16288
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 14176 4527 15200
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 13088 4527 14112
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 12000 4527 13024
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 10912 4527 11936
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 9824 4527 10848
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 8736 4527 9760
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 7648 4527 8672
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 6560 4527 7584
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 5472 4527 6496
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 4384 4527 5408
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 3296 4527 4320
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 2208 4527 3232
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2128 4527 2144
rect 5839 41920 6159 42944
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 40832 6159 41856
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 39744 6159 40768
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 38656 6159 39680
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 37568 6159 38592
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 36480 6159 37504
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 35392 6159 36416
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 34304 6159 35328
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 33216 6159 34240
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 32128 6159 33152
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 31040 6159 32064
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 29952 6159 30976
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 28864 6159 29888
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 27776 6159 28800
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 26688 6159 27712
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 25600 6159 26624
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 24512 6159 25536
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 23424 6159 24448
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 22336 6159 23360
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 21248 6159 22272
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 20160 6159 21184
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 19072 6159 20096
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 17984 6159 19008
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 16896 6159 17920
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 15808 6159 16832
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 14720 6159 15744
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 13632 6159 14656
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 12544 6159 13568
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 11456 6159 12480
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 10368 6159 11392
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 9280 6159 10304
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 8192 6159 9216
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 7104 6159 8128
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 6016 6159 7040
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 4928 6159 5952
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 3840 6159 4864
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 2752 6159 3776
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2128 6159 2688
rect 7471 43552 7791 44576
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 42464 7791 43488
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 41376 7791 42400
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 7471 40288 7791 41312
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 39200 7791 40224
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 38112 7791 39136
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 37024 7791 38048
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 35936 7791 36960
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 34848 7791 35872
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 33760 7791 34784
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 32672 7791 33696
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 31584 7791 32608
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 30496 7791 31520
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 29408 7791 30432
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 28320 7791 29344
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 27232 7791 28256
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 26144 7791 27168
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 25056 7791 26080
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 23968 7791 24992
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 22880 7791 23904
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 21792 7791 22816
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 20704 7791 21728
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 19616 7791 20640
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 18528 7791 19552
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 17440 7791 18464
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 16352 7791 17376
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 15264 7791 16288
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 14176 7791 15200
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 13088 7791 14112
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 12000 7791 13024
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 10912 7791 11936
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 9824 7791 10848
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 8736 7791 9760
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 7648 7791 8672
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 6560 7791 7584
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 5472 7791 6496
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 4384 7791 5408
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 3296 7791 4320
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 2208 7791 3232
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2128 7791 2144
rect 9103 77824 9423 77840
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 76736 9423 77760
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 75648 9423 76672
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 74560 9423 75584
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 73472 9423 74496
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 72384 9423 73408
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 71296 9423 72320
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 70208 9423 71232
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 69120 9423 70144
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 68032 9423 69056
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 66944 9423 67968
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 65856 9423 66880
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 64768 9423 65792
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 63680 9423 64704
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 62592 9423 63616
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 61504 9423 62528
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 60416 9423 61440
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 59328 9423 60352
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 58240 9423 59264
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 57152 9423 58176
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 56064 9423 57088
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 54976 9423 56000
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 53888 9423 54912
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 52800 9423 53824
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 51712 9423 52736
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 50624 9423 51648
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 49536 9423 50560
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 48448 9423 49472
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 47360 9423 48384
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 46272 9423 47296
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 45184 9423 46208
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 44096 9423 45120
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 43008 9423 44032
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 41920 9423 42944
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 40832 9423 41856
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 39744 9423 40768
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 38656 9423 39680
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 37568 9423 38592
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 36480 9423 37504
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 35392 9423 36416
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 34304 9423 35328
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 33216 9423 34240
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 32128 9423 33152
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 31040 9423 32064
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 29952 9423 30976
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 28864 9423 29888
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 27776 9423 28800
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 26688 9423 27712
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 25600 9423 26624
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 24512 9423 25536
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 23424 9423 24448
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 22336 9423 23360
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 21248 9423 22272
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 20160 9423 21184
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 19072 9423 20096
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 17984 9423 19008
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 16896 9423 17920
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 15808 9423 16832
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 14720 9423 15744
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 13632 9423 14656
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 12544 9423 13568
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 11456 9423 12480
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 10368 9423 11392
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 9280 9423 10304
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 8192 9423 9216
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 7104 9423 8128
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 6016 9423 7040
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 4928 9423 5952
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 3840 9423 4864
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 2752 9423 3776
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2128 9423 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1635444444
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1635444444
transform -1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1635444444
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1635444444
transform 1 0 2392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1635444444
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _261_
timestamp 1635444444
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1635444444
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1635444444
transform 1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1635444444
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1635444444
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4324 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1635444444
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1635444444
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39
timestamp 1635444444
transform 1 0 4692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46
timestamp 1635444444
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1635444444
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1635444444
transform 1 0 5060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1635444444
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1635444444
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1635444444
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1635444444
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1635444444
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1635444444
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1635444444
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1635444444
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1635444444
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1635444444
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1635444444
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1635444444
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1635444444
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1635444444
transform 1 0 1380 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _224_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2760 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1635444444
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1635444444
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1635444444
transform 1 0 4048 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1635444444
transform 1 0 5152 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1635444444
transform 1 0 6256 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1635444444
transform 1 0 7360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1635444444
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1635444444
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1635444444
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1635444444
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1635444444
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1635444444
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _223_
timestamp 1635444444
transform -1 0 2852 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1635444444
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 1635444444
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_33
timestamp 1635444444
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _181_
timestamp 1635444444
transform -1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1635444444
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1635444444
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1635444444
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1635444444
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1635444444
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1635444444
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1635444444
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1635444444
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _186_
timestamp 1635444444
transform -1 0 3036 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1635444444
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1635444444
transform 1 0 4048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1635444444
transform 1 0 5152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1635444444
transform 1 0 6256 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1635444444
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1635444444
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1635444444
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1635444444
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1635444444
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1635444444
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1635444444
transform -1 0 2392 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _262_
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1635444444
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_21
timestamp 1635444444
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _183_
timestamp 1635444444
transform -1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _185_
timestamp 1635444444
transform -1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1635444444
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_35
timestamp 1635444444
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _187_
timestamp 1635444444
transform -1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1635444444
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635444444
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1635444444
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1635444444
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1635444444
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1635444444
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1635444444
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_12
timestamp 1635444444
transform 1 0 2208 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_6
timestamp 1635444444
transform 1 0 1656 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 1635444444
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1635444444
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1635444444
transform -1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_16
timestamp 1635444444
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1635444444
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_20
timestamp 1635444444
transform 1 0 2944 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1635444444
transform -1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1635444444
transform -1 0 2944 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1635444444
transform -1 0 3588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1635444444
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1635444444
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1635444444
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1635444444
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1635444444
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1635444444
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1635444444
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1635444444
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1635444444
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1635444444
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1635444444
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1635444444
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1635444444
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1635444444
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1635444444
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1635444444
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_7
timestamp 1635444444
transform 1 0 1748 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input97
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_15
timestamp 1635444444
transform 1 0 2484 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1635444444
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _238_
timestamp 1635444444
transform -1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1635444444
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1635444444
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1635444444
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1635444444
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1635444444
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1635444444
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1635444444
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1635444444
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1635444444
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 1635444444
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1635444444
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _188_
timestamp 1635444444
transform -1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1635444444
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _189_
timestamp 1635444444
transform -1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input98
timestamp 1635444444
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1635444444
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1635444444
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1635444444
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1635444444
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1635444444
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1635444444
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1635444444
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1635444444
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1635444444
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_10_13
timestamp 1635444444
transform 1 0 2300 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_20
timestamp 1635444444
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1635444444
transform -1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1635444444
transform 1 0 4048 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1635444444
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1635444444
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1635444444
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1635444444
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1635444444
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1635444444
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1635444444
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _263_
timestamp 1635444444
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _266_
timestamp 1635444444
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_15
timestamp 1635444444
transform 1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1635444444
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1635444444
transform -1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_29
timestamp 1635444444
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1635444444
transform -1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_41
timestamp 1635444444
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1635444444
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1635444444
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1635444444
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_93
timestamp 1635444444
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1635444444
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1635444444
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1635444444
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1635444444
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _264_
timestamp 1635444444
transform -1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_17
timestamp 1635444444
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1635444444
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _265_
timestamp 1635444444
transform -1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1635444444
transform -1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1635444444
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1635444444
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1635444444
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1635444444
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1635444444
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1635444444
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _247_
timestamp 1635444444
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp 1635444444
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1635444444
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1635444444
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1635444444
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1635444444
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_22
timestamp 1635444444
transform 1 0 3128 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1635444444
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1635444444
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _241_
timestamp 1635444444
transform -1 0 2944 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_34
timestamp 1635444444
transform 1 0 4232 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1635444444
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1635444444
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1635444444
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1635444444
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1635444444
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1635444444
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1635444444
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_81
timestamp 1635444444
transform 1 0 8556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_87
timestamp 1635444444
transform 1 0 9108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1635444444
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _249_
timestamp 1635444444
transform -1 0 9476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _250_
timestamp 1635444444
transform -1 0 9568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 1635444444
transform 1 0 9476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1635444444
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1635444444
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1635444444
transform 1 0 10212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1635444444
transform 1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1635444444
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1635444444
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _225_
timestamp 1635444444
transform 1 0 2668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1635444444
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1635444444
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1635444444
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1635444444
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1635444444
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1635444444
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1635444444
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1635444444
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1635444444
transform 1 0 1380 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1635444444
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_20
timestamp 1635444444
transform 1 0 2944 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _242_
timestamp 1635444444
transform -1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1635444444
transform 1 0 4048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1635444444
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1635444444
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1635444444
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1635444444
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1635444444
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1635444444
transform 1 0 9660 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1635444444
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1635444444
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1635444444
transform 1 0 1380 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1635444444
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_21
timestamp 1635444444
transform 1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1635444444
transform -1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _267_
timestamp 1635444444
transform -1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_28
timestamp 1635444444
transform 1 0 3680 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_35
timestamp 1635444444
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _245_
timestamp 1635444444
transform -1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1635444444
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1635444444
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1635444444
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1635444444
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1635444444
transform 1 0 10396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_93
timestamp 1635444444
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1635444444
transform 1 0 1380 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1635444444
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1635444444
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _268_
timestamp 1635444444
transform -1 0 3036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1635444444
transform 1 0 4048 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _246_
timestamp 1635444444
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1635444444
transform 1 0 5152 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1635444444
transform 1 0 6256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1635444444
transform 1 0 7360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1635444444
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1635444444
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1635444444
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1635444444
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1635444444
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1635444444
transform 1 0 1380 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1635444444
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_21
timestamp 1635444444
transform 1 0 3036 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1635444444
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1635444444
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _269_
timestamp 1635444444
transform -1 0 3036 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_33
timestamp 1635444444
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1635444444
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1635444444
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1635444444
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1635444444
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1635444444
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1635444444
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1635444444
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1635444444
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1635444444
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1635444444
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1635444444
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1635444444
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_97
timestamp 1635444444
transform 1 0 10028 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1635444444
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_11
timestamp 1635444444
transform 1 0 2116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1635444444
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1635444444
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_20
timestamp 1635444444
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_32
timestamp 1635444444
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1635444444
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1635444444
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_81
timestamp 1635444444
transform 1 0 8556 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 1635444444
transform 1 0 9108 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _251_
timestamp 1635444444
transform -1 0 9476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_91
timestamp 1635444444
transform 1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1635444444
transform 1 0 10212 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1635444444
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_9
timestamp 1635444444
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_16
timestamp 1635444444
transform 1 0 2576 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1635444444
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1635444444
transform 1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1635444444
transform 1 0 2944 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1635444444
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1635444444
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1635444444
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1635444444
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1635444444
transform 1 0 7360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1635444444
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1635444444
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1635444444
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1635444444
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_11
timestamp 1635444444
transform 1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1635444444
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _067_
timestamp 1635444444
transform 1 0 1656 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_23_21
timestamp 1635444444
transform 1 0 3036 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_1  _068_
timestamp 1635444444
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_33
timestamp 1635444444
transform 1 0 4140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_45
timestamp 1635444444
transform 1 0 5244 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1635444444
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1635444444
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1635444444
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1635444444
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1635444444
transform 1 0 10212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1635444444
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1635444444
transform 1 0 1656 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _061_
timestamp 1635444444
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1635444444
transform 1 0 2024 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_13
timestamp 1635444444
transform 1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1635444444
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1635444444
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1635444444
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1635444444
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1635444444
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1635444444
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1635444444
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1635444444
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1635444444
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1635444444
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1635444444
transform 1 0 2024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1635444444
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _063_
timestamp 1635444444
transform 1 0 1472 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_19
timestamp 1635444444
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__nand4_1  _066_
timestamp 1635444444
transform 1 0 2392 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_25_31
timestamp 1635444444
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_43
timestamp 1635444444
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1635444444
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1635444444
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1635444444
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1635444444
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1635444444
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1635444444
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1635444444
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1635444444
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1635444444
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1635444444
transform -1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1635444444
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1635444444
transform 1 0 2024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1635444444
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1635444444
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_20
timestamp 1635444444
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1635444444
transform 1 0 2668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1635444444
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1635444444
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1635444444
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1635444444
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1635444444
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1635444444
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1635444444
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1635444444
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1635444444
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1635444444
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1635444444
transform -1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_91
timestamp 1635444444
transform 1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1635444444
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_93
timestamp 1635444444
transform 1 0 9660 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1635444444
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _253_
timestamp 1635444444
transform 1 0 9936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1635444444
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_11
timestamp 1635444444
transform 1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1635444444
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1635444444
transform 1 0 1748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1635444444
transform -1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 1635444444
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1635444444
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1635444444
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1635444444
transform 1 0 4048 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1635444444
transform 1 0 5152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1635444444
transform 1 0 6256 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1635444444
transform 1 0 7360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1635444444
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1635444444
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_99
timestamp 1635444444
transform 1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1635444444
transform 1 0 9844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1635444444
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_8
timestamp 1635444444
transform 1 0 1840 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1635444444
transform -1 0 1840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_19
timestamp 1635444444
transform 1 0 2852 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2852 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1635444444
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1635444444
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1635444444
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_50
timestamp 1635444444
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1635444444
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_81
timestamp 1635444444
transform 1 0 8556 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_87
timestamp 1635444444
transform 1 0 9108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1635444444
transform -1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_91
timestamp 1635444444
transform 1 0 9476 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_99
timestamp 1635444444
transform 1 0 10212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1635444444
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_8
timestamp 1635444444
transform 1 0 1840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _070_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2208 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__clkinv_2  _079_
timestamp 1635444444
transform -1 0 1840 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1635444444
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1635444444
transform 1 0 4048 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1635444444
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1635444444
transform 1 0 6256 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1635444444
transform 1 0 7360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1635444444
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _255_
timestamp 1635444444
transform -1 0 9476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1635444444
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1635444444
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1635444444
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1635444444
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1635444444
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _081_
timestamp 1635444444
transform -1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_16
timestamp 1635444444
transform 1 0 2576 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1635444444
transform -1 0 2576 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_28
timestamp 1635444444
transform 1 0 3680 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_40
timestamp 1635444444
transform 1 0 4784 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1635444444
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1635444444
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1635444444
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1635444444
transform 1 0 10488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_93
timestamp 1635444444
transform 1 0 9660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1635444444
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _257_
timestamp 1635444444
transform 1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_9
timestamp 1635444444
transform 1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _083_
timestamp 1635444444
transform -1 0 1932 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1635444444
transform 1 0 2576 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1635444444
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1635444444
transform 1 0 2300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1635444444
transform 1 0 2944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1635444444
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1635444444
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1635444444
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1635444444
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1635444444
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1635444444
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1635444444
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1635444444
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1635444444
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1635444444
transform -1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1635444444
transform 1 0 1380 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1635444444
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1635444444
transform -1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_7
timestamp 1635444444
transform 1 0 1748 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_7
timestamp 1635444444
transform 1 0 1748 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _089_
timestamp 1635444444
transform -1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_11
timestamp 1635444444
transform 1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_18
timestamp 1635444444
transform 1 0 2760 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_25
timestamp 1635444444
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 1635444444
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_23
timestamp 1635444444
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _091_
timestamp 1635444444
transform 1 0 2852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1635444444
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1635444444
transform 1 0 3128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_37
timestamp 1635444444
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1635444444
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1635444444
transform 1 0 4048 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1635444444
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1635444444
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1635444444
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1635444444
transform 1 0 6256 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1635444444
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1635444444
transform 1 0 7360 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_81
timestamp 1635444444
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1635444444
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1635444444
transform 1 0 9660 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1635444444
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_102
timestamp 1635444444
transform 1 0 10488 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1635444444
transform 1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_98
timestamp 1635444444
transform 1 0 10120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1635444444
transform 1 0 9844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1635444444
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_6
timestamp 1635444444
transform 1 0 1656 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1635444444
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_14
timestamp 1635444444
transform 1 0 2392 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_21
timestamp 1635444444
transform 1 0 3036 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__or2b_1  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2484 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_33
timestamp 1635444444
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_45
timestamp 1635444444
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1635444444
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1635444444
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1635444444
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_93
timestamp 1635444444
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_99
timestamp 1635444444
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1635444444
transform 1 0 9844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_7
timestamp 1635444444
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2576 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1635444444
transform -1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_16
timestamp 1635444444
transform 1 0 2576 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_23
timestamp 1635444444
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1635444444
transform 1 0 2944 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1635444444
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1635444444
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1635444444
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1635444444
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1635444444
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1635444444
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _259_
timestamp 1635444444
transform -1 0 9476 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_91
timestamp 1635444444
transform 1 0 9476 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1635444444
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_6
timestamp 1635444444
transform 1 0 1656 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1635444444
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _071_
timestamp 1635444444
transform 1 0 2392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_26
timestamp 1635444444
transform 1 0 3496 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_33
timestamp 1635444444
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1635444444
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1635444444
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1635444444
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1635444444
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1635444444
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1635444444
transform 1 0 9660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1635444444
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1635444444
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_11
timestamp 1635444444
transform 1 0 2116 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1635444444
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _074_
timestamp 1635444444
transform 1 0 1656 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_38_17
timestamp 1635444444
transform 1 0 2668 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1635444444
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _137_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2760 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1635444444
transform 1 0 4048 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _190_
timestamp 1635444444
transform -1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1635444444
transform 1 0 5152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1635444444
transform 1 0 6256 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1635444444
transform 1 0 7360 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1635444444
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp 1635444444
transform -1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_92
timestamp 1635444444
transform 1 0 9568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1635444444
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_6
timestamp 1635444444
transform 1 0 1656 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1635444444
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_9
timestamp 1635444444
transform 1 0 1932 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _076_
timestamp 1635444444
transform 1 0 2024 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _103_
timestamp 1635444444
transform -1 0 1932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1635444444
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_15
timestamp 1635444444
transform 1 0 2484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_24
timestamp 1635444444
transform 1 0 3312 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_20
timestamp 1635444444
transform 1 0 2944 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _191_
timestamp 1635444444
transform -1 0 2944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _226_
timestamp 1635444444
transform -1 0 3312 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_39_31
timestamp 1635444444
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1635444444
transform 1 0 4048 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _192_
timestamp 1635444444
transform -1 0 3956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_43
timestamp 1635444444
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1635444444
transform 1 0 5152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1635444444
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1635444444
transform 1 0 6256 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1635444444
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1635444444
transform 1 0 7360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1635444444
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1635444444
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1635444444
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_93
timestamp 1635444444
transform 1 0 9660 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1635444444
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_97
timestamp 1635444444
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1635444444
transform 1 0 9844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_10
timestamp 1635444444
transform 1 0 2024 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_6
timestamp 1635444444
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1635444444
transform 1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1635444444
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_14
timestamp 1635444444
transform 1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_21
timestamp 1635444444
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1635444444
transform 1 0 2760 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_33
timestamp 1635444444
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1635444444
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1635444444
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1635444444
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_93
timestamp 1635444444
transform 1 0 9660 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1635444444
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _232_
timestamp 1635444444
transform 1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_10
timestamp 1635444444
transform 1 0 2024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _108_
timestamp 1635444444
transform -1 0 2024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_17
timestamp 1635444444
transform 1 0 2668 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_25
timestamp 1635444444
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1635444444
transform 1 0 2392 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1635444444
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1635444444
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1635444444
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_93
timestamp 1635444444
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1635444444
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _233_
timestamp 1635444444
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_6
timestamp 1635444444
transform 1 0 1656 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1635444444
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1635444444
transform -1 0 2300 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_13
timestamp 1635444444
transform 1 0 2300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_20
timestamp 1635444444
transform 1 0 2944 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1635444444
transform 1 0 2668 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_32
timestamp 1635444444
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_44
timestamp 1635444444
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1635444444
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1635444444
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_101
timestamp 1635444444
transform 1 0 10396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1635444444
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_7
timestamp 1635444444
transform 1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _110_
timestamp 1635444444
transform 1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _112_
timestamp 1635444444
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_15
timestamp 1635444444
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1635444444
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1635444444
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1635444444
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1635444444
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1635444444
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1635444444
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1635444444
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1635444444
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_93
timestamp 1635444444
transform 1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_99
timestamp 1635444444
transform 1 0 10212 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _234_
timestamp 1635444444
transform 1 0 9936 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1635444444
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1635444444
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _118_
timestamp 1635444444
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_16
timestamp 1635444444
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_23
timestamp 1635444444
transform 1 0 3220 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1635444444
transform -1 0 2576 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1635444444
transform 1 0 2944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_35
timestamp 1635444444
transform 1 0 4324 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_47
timestamp 1635444444
transform 1 0 5428 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1635444444
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1635444444
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1635444444
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_101
timestamp 1635444444
transform 1 0 10396 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_93
timestamp 1635444444
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1635444444
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_3
timestamp 1635444444
transform 1 0 1380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_8
timestamp 1635444444
transform 1 0 1840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _116_
timestamp 1635444444
transform 1 0 2024 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _120_
timestamp 1635444444
transform -1 0 1840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1635444444
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1635444444
transform 1 0 2208 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_14
timestamp 1635444444
transform 1 0 2392 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1635444444
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1635444444
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1635444444
transform 1 0 2760 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1635444444
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_29
timestamp 1635444444
transform 1 0 3772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1635444444
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4140 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1635444444
transform 1 0 5152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1635444444
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1635444444
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1635444444
transform 1 0 6256 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1635444444
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1635444444
transform 1 0 7360 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1635444444
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1635444444
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1635444444
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1635444444
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_101
timestamp 1635444444
transform 1 0 10396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_93
timestamp 1635444444
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _229_
timestamp 1635444444
transform -1 0 10212 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_3
timestamp 1635444444
transform 1 0 1380 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_8
timestamp 1635444444
transform 1 0 1840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1635444444
transform -1 0 2484 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _122_
timestamp 1635444444
transform -1 0 1840 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_15
timestamp 1635444444
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_22
timestamp 1635444444
transform 1 0 3128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1635444444
transform -1 0 3128 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1635444444
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1635444444
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1635444444
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1635444444
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1635444444
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1635444444
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_93
timestamp 1635444444
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_99
timestamp 1635444444
transform 1 0 10212 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _230_
timestamp 1635444444
transform -1 0 10212 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_6
timestamp 1635444444
transform 1 0 1656 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _228_
timestamp 1635444444
transform -1 0 2668 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1635444444
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_17
timestamp 1635444444
transform 1 0 2668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_24
timestamp 1635444444
transform 1 0 3312 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1635444444
transform 1 0 3036 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_36
timestamp 1635444444
transform 1 0 4416 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1635444444
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1635444444
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_101
timestamp 1635444444
transform 1 0 10396 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_93
timestamp 1635444444
transform 1 0 9660 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_3
timestamp 1635444444
transform 1 0 1380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_8
timestamp 1635444444
transform 1 0 1840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _124_
timestamp 1635444444
transform 1 0 1472 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _227_
timestamp 1635444444
transform -1 0 2668 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_50_17
timestamp 1635444444
transform 1 0 2668 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1635444444
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _193_
timestamp 1635444444
transform -1 0 3312 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1635444444
transform 1 0 4048 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1635444444
transform 1 0 5152 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_56
timestamp 1635444444
transform 1 0 6256 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_68
timestamp 1635444444
transform 1 0 7360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1635444444
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_97
timestamp 1635444444
transform 1 0 10028 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_7
timestamp 1635444444
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _078_
timestamp 1635444444
transform -1 0 2576 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1635444444
transform -1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_16
timestamp 1635444444
transform 1 0 2576 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_24
timestamp 1635444444
transform 1 0 3312 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _126_
timestamp 1635444444
transform 1 0 2944 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_31
timestamp 1635444444
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1635444444
transform 1 0 3680 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_43
timestamp 1635444444
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1635444444
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1635444444
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1635444444
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_93
timestamp 1635444444
transform 1 0 9660 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_99
timestamp 1635444444
transform 1 0 10212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _235_
timestamp 1635444444
transform 1 0 9936 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_3
timestamp 1635444444
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_9
timestamp 1635444444
transform 1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _128_
timestamp 1635444444
transform -1 0 2300 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _130_
timestamp 1635444444
transform -1 0 1932 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_13
timestamp 1635444444
transform 1 0 2300 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_20
timestamp 1635444444
transform 1 0 2944 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_17
timestamp 1635444444
transform 1 0 2668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1635444444
transform -1 0 2944 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _132_
timestamp 1635444444
transform -1 0 2668 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1635444444
transform 1 0 4048 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_29
timestamp 1635444444
transform 1 0 3772 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1635444444
transform 1 0 5152 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_41
timestamp 1635444444
transform 1 0 4876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_56
timestamp 1635444444
transform 1 0 6256 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1635444444
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1635444444
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_68
timestamp 1635444444
transform 1 0 7360 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1635444444
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1635444444
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_85
timestamp 1635444444
transform 1 0 8924 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1635444444
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _236_
timestamp 1635444444
transform 1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_91
timestamp 1635444444
transform 1 0 9476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1635444444
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1635444444
transform 1 0 9660 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1635444444
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1635444444
transform 1 0 9844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1635444444
transform 1 0 9844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_11
timestamp 1635444444
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _134_
timestamp 1635444444
transform -1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 1635444444
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1635444444
transform 1 0 2484 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1635444444
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1635444444
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1635444444
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1635444444
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1635444444
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1635444444
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1635444444
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1635444444
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1635444444
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1635444444
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_7
timestamp 1635444444
transform 1 0 1748 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1635444444
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_15
timestamp 1635444444
transform 1 0 2484 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_21
timestamp 1635444444
transform 1 0 3036 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _194_
timestamp 1635444444
transform -1 0 3036 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_33
timestamp 1635444444
transform 1 0 4140 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_45
timestamp 1635444444
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_53
timestamp 1635444444
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1635444444
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1635444444
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1635444444
transform 1 0 10396 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_93
timestamp 1635444444
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1635444444
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1635444444
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1635444444
transform 1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_15
timestamp 1635444444
transform 1 0 2484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_22
timestamp 1635444444
transform 1 0 3128 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _195_
timestamp 1635444444
transform -1 0 3128 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1635444444
transform 1 0 4048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1635444444
transform -1 0 4048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1635444444
transform 1 0 5152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1635444444
transform 1 0 6256 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1635444444
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1635444444
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_93
timestamp 1635444444
transform 1 0 9660 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_99
timestamp 1635444444
transform 1 0 10212 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1635444444
transform 1 0 9844 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1635444444
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1635444444
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1635444444
transform 1 0 2116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_15
timestamp 1635444444
transform 1 0 2484 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_22
timestamp 1635444444
transform 1 0 3128 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1635444444
transform 1 0 2852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_34
timestamp 1635444444
transform 1 0 4232 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_46
timestamp 1635444444
transform 1 0 5336 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1635444444
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1635444444
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1635444444
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_93
timestamp 1635444444
transform 1 0 9660 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_99
timestamp 1635444444
transform 1 0 10212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1635444444
transform 1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_7
timestamp 1635444444
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1635444444
transform -1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1635444444
transform 1 0 2116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_15
timestamp 1635444444
transform 1 0 2484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_22
timestamp 1635444444
transform 1 0 3128 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _198_
timestamp 1635444444
transform -1 0 3128 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1635444444
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1635444444
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1635444444
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1635444444
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1635444444
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1635444444
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_97
timestamp 1635444444
transform 1 0 10028 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_3
timestamp 1635444444
transform 1 0 1380 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_9
timestamp 1635444444
transform 1 0 1932 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_3
timestamp 1635444444
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_7
timestamp 1635444444
transform 1 0 1748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _082_
timestamp 1635444444
transform 1 0 1840 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _088_
timestamp 1635444444
transform 1 0 1472 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_59_17
timestamp 1635444444
transform 1 0 2668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_25
timestamp 1635444444
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_13
timestamp 1635444444
transform 1 0 2300 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_22
timestamp 1635444444
transform 1 0 3128 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _086_
timestamp 1635444444
transform -1 0 3128 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1635444444
transform -1 0 2668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1635444444
transform 1 0 3036 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_37
timestamp 1635444444
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1635444444
transform 1 0 4048 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _197_
timestamp 1635444444
transform -1 0 4048 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1635444444
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1635444444
transform 1 0 5152 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1635444444
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1635444444
transform 1 0 6256 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1635444444
transform 1 0 7360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1635444444
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1635444444
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_93
timestamp 1635444444
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_99
timestamp 1635444444
transform 1 0 10212 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1635444444
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1635444444
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1635444444
transform 1 0 9844 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1635444444
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1635444444
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _080_
timestamp 1635444444
transform -1 0 2484 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_61_15
timestamp 1635444444
transform 1 0 2484 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_23
timestamp 1635444444
transform 1 0 3220 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1635444444
transform 1 0 2852 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_35
timestamp 1635444444
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1635444444
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1635444444
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1635444444
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1635444444
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_101
timestamp 1635444444
transform 1 0 10396 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_93
timestamp 1635444444
transform 1 0 9660 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_12
timestamp 1635444444
transform 1 0 2208 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1635444444
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _084_
timestamp 1635444444
transform -1 0 2208 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_62_20
timestamp 1635444444
transform 1 0 2944 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1635444444
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _199_
timestamp 1635444444
transform -1 0 3312 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1635444444
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1635444444
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1635444444
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1635444444
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1635444444
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1635444444
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1635444444
transform 1 0 9660 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1635444444
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1635444444
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1635444444
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1635444444
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1635444444
transform 1 0 2116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1635444444
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_23
timestamp 1635444444
transform 1 0 3220 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1635444444
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_35
timestamp 1635444444
transform 1 0 4324 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1635444444
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1635444444
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1635444444
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_93
timestamp 1635444444
transform 1 0 9660 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_99
timestamp 1635444444
transform 1 0 10212 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1635444444
transform 1 0 9844 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_3
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_9
timestamp 1635444444
transform 1 0 1932 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _094_
timestamp 1635444444
transform 1 0 1472 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_64_18
timestamp 1635444444
transform 1 0 2760 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _202_
timestamp 1635444444
transform -1 0 2760 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_26
timestamp 1635444444
transform 1 0 3496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1635444444
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1635444444
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1635444444
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1635444444
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1635444444
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1635444444
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1635444444
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1635444444
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_99
timestamp 1635444444
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1635444444
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_7
timestamp 1635444444
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _092_
timestamp 1635444444
transform -1 0 2576 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1635444444
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_16
timestamp 1635444444
transform 1 0 2576 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_25
timestamp 1635444444
transform 1 0 3404 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _096_
timestamp 1635444444
transform -1 0 3404 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_65_37
timestamp 1635444444
transform 1 0 4508 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_49
timestamp 1635444444
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1635444444
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1635444444
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1635444444
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_101
timestamp 1635444444
transform 1 0 10396 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_93
timestamp 1635444444
transform 1 0 9660 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_7
timestamp 1635444444
transform 1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_11
timestamp 1635444444
transform 1 0 2116 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1635444444
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _090_
timestamp 1635444444
transform -1 0 2576 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _270_
timestamp 1635444444
transform 1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1635444444
transform -1 0 1748 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_16
timestamp 1635444444
transform 1 0 2576 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_23
timestamp 1635444444
transform 1 0 3220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_19
timestamp 1635444444
transform 1 0 2852 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _203_
timestamp 1635444444
transform -1 0 3220 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1635444444
transform -1 0 2852 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1635444444
transform 1 0 3220 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1635444444
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1635444444
transform 1 0 4048 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_27
timestamp 1635444444
transform 1 0 3588 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_34
timestamp 1635444444
transform 1 0 4232 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1635444444
transform -1 0 4048 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _204_
timestamp 1635444444
transform -1 0 4232 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1635444444
transform 1 0 5152 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_46
timestamp 1635444444
transform 1 0 5336 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1635444444
transform 1 0 6256 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1635444444
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1635444444
transform 1 0 7360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1635444444
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1635444444
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_85
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1635444444
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_93
timestamp 1635444444
transform 1 0 9660 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_99
timestamp 1635444444
transform 1 0 10212 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_93
timestamp 1635444444
transform 1 0 9660 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_99
timestamp 1635444444
transform 1 0 10212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1635444444
transform 1 0 9844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1635444444
transform 1 0 9844 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_10
timestamp 1635444444
transform 1 0 2024 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1635444444
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _098_
timestamp 1635444444
transform -1 0 2024 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_68_18
timestamp 1635444444
transform 1 0 2760 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1635444444
transform 1 0 2392 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_26
timestamp 1635444444
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1635444444
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1635444444
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1635444444
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1635444444
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1635444444
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1635444444
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_97
timestamp 1635444444
transform 1 0 10028 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_7
timestamp 1635444444
transform 1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _102_
timestamp 1635444444
transform 1 0 2116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1635444444
transform -1 0 1748 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_14
timestamp 1635444444
transform 1 0 2392 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_18
timestamp 1635444444
transform 1 0 2760 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_22
timestamp 1635444444
transform 1 0 3128 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _205_
timestamp 1635444444
transform -1 0 3128 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_34
timestamp 1635444444
transform 1 0 4232 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_46
timestamp 1635444444
transform 1 0 5336 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_54
timestamp 1635444444
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1635444444
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1635444444
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_93
timestamp 1635444444
transform 1 0 9660 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_99
timestamp 1635444444
transform 1 0 10212 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1635444444
transform 1 0 9844 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_7
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _100_
timestamp 1635444444
transform 1 0 2116 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1635444444
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_14
timestamp 1635444444
transform 1 0 2392 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_26
timestamp 1635444444
transform 1 0 3496 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1635444444
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1635444444
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1635444444
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1635444444
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1635444444
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_85
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_93
timestamp 1635444444
transform 1 0 9660 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_99
timestamp 1635444444
transform 1 0 10212 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1635444444
transform 1 0 9844 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_7
timestamp 1635444444
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1635444444
transform -1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1635444444
transform -1 0 2484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_15
timestamp 1635444444
transform 1 0 2484 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_23
timestamp 1635444444
transform 1 0 3220 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1635444444
transform 1 0 2852 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_35
timestamp 1635444444
transform 1 0 4324 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_47
timestamp 1635444444
transform 1 0 5428 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1635444444
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1635444444
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_93
timestamp 1635444444
transform 1 0 9660 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1635444444
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1635444444
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_3
timestamp 1635444444
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _113_
timestamp 1635444444
transform -1 0 2392 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1635444444
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1635444444
transform -1 0 2484 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_14
timestamp 1635444444
transform 1 0 2392 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1635444444
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_73_15
timestamp 1635444444
transform 1 0 2484 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_21
timestamp 1635444444
transform 1 0 3036 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_25
timestamp 1635444444
transform 1 0 3404 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _206_
timestamp 1635444444
transform -1 0 3036 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _208_
timestamp 1635444444
transform -1 0 3404 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1635444444
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_37
timestamp 1635444444
transform 1 0 4508 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1635444444
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_49
timestamp 1635444444
transform 1 0 5612 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1635444444
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1635444444
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1635444444
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1635444444
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1635444444
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1635444444
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1635444444
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_97
timestamp 1635444444
transform 1 0 10028 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_93
timestamp 1635444444
transform 1 0 9660 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_99
timestamp 1635444444
transform 1 0 10212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1635444444
transform 1 0 9844 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_6
timestamp 1635444444
transform 1 0 1656 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _107_
timestamp 1635444444
transform -1 0 1656 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _115_
timestamp 1635444444
transform -1 0 2484 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_74_15
timestamp 1635444444
transform 1 0 2484 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_23
timestamp 1635444444
transform 1 0 3220 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1635444444
transform 1 0 2852 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635444444
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1635444444
transform 1 0 4048 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _212_
timestamp 1635444444
transform -1 0 4048 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1635444444
transform 1 0 5152 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_56
timestamp 1635444444
transform 1 0 6256 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1635444444
transform 1 0 7360 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_80
timestamp 1635444444
transform 1 0 8464 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_93
timestamp 1635444444
transform 1 0 9660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_99
timestamp 1635444444
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1635444444
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_11
timestamp 1635444444
transform 1 0 2116 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_3
timestamp 1635444444
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _119_
timestamp 1635444444
transform -1 0 2116 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_75_19
timestamp 1635444444
transform 1 0 2852 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _105_
timestamp 1635444444
transform 1 0 3220 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1635444444
transform 1 0 2484 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_26
timestamp 1635444444
transform 1 0 3496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_33
timestamp 1635444444
transform 1 0 4140 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _209_
timestamp 1635444444
transform -1 0 4140 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1635444444
transform -1 0 4784 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_40
timestamp 1635444444
transform 1 0 4784 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1635444444
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1635444444
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1635444444
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_101
timestamp 1635444444
transform 1 0 10396 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_93
timestamp 1635444444
transform 1 0 9660 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_76_3
timestamp 1635444444
transform 1 0 1380 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_9
timestamp 1635444444
transform 1 0 1932 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _121_
timestamp 1635444444
transform -1 0 1932 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_76_17
timestamp 1635444444
transform 1 0 2668 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1635444444
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _207_
timestamp 1635444444
transform -1 0 3312 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1635444444
transform -1 0 2668 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1635444444
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1635444444
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1635444444
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1635444444
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1635444444
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_93
timestamp 1635444444
transform 1 0 9660 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_99
timestamp 1635444444
transform 1 0 10212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1635444444
transform 1 0 9844 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_77_7
timestamp 1635444444
transform 1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1635444444
transform -1 0 1748 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1635444444
transform 1 0 2116 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_15
timestamp 1635444444
transform 1 0 2484 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_23
timestamp 1635444444
transform 1 0 3220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1635444444
transform -1 0 3220 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_30
timestamp 1635444444
transform 1 0 3864 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _210_
timestamp 1635444444
transform -1 0 3864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_42
timestamp 1635444444
transform 1 0 4968 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_54
timestamp 1635444444
transform 1 0 6072 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1635444444
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1635444444
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_93
timestamp 1635444444
transform 1 0 9660 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_99
timestamp 1635444444
transform 1 0 10212 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1635444444
transform 1 0 9844 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_11
timestamp 1635444444
transform 1 0 2116 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_3
timestamp 1635444444
transform 1 0 1380 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _123_
timestamp 1635444444
transform 1 0 1656 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_78_19
timestamp 1635444444
transform 1 0 2852 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1635444444
transform 1 0 2484 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1635444444
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1635444444
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1635444444
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1635444444
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1635444444
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1635444444
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1635444444
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_93
timestamp 1635444444
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1635444444
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1635444444
transform 1 0 9844 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_7
timestamp 1635444444
transform 1 0 1748 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1635444444
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _271_
timestamp 1635444444
transform 1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1635444444
transform -1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1635444444
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_14
timestamp 1635444444
transform 1 0 2392 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_19
timestamp 1635444444
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_26
timestamp 1635444444
transform 1 0 3496 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_38
timestamp 1635444444
transform 1 0 4600 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1635444444
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1635444444
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_79_50
timestamp 1635444444
transform 1 0 5704 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1635444444
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1635444444
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1635444444
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1635444444
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1635444444
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1635444444
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1635444444
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_85
timestamp 1635444444
transform 1 0 8924 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_101
timestamp 1635444444
transform 1 0 10396 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_93
timestamp 1635444444
transform 1 0 9660 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_93
timestamp 1635444444
transform 1 0 9660 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_99
timestamp 1635444444
transform 1 0 10212 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1635444444
transform 1 0 9844 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1635444444
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_81_7
timestamp 1635444444
transform 1 0 1748 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1635444444
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1635444444
transform -1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_18
timestamp 1635444444
transform 1 0 2760 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _215_
timestamp 1635444444
transform -1 0 2760 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_30
timestamp 1635444444
transform 1 0 3864 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_42
timestamp 1635444444
transform 1 0 4968 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1635444444
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1635444444
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1635444444
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1635444444
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_93
timestamp 1635444444
transform 1 0 9660 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1635444444
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1635444444
transform 1 0 9844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1635444444
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_11
timestamp 1635444444
transform 1 0 2116 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_7
timestamp 1635444444
transform 1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1635444444
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _117_
timestamp 1635444444
transform -1 0 2484 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1635444444
transform -1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_15
timestamp 1635444444
transform 1 0 2484 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_22
timestamp 1635444444
transform 1 0 3128 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _214_
timestamp 1635444444
transform -1 0 3128 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1635444444
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1635444444
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1635444444
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1635444444
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1635444444
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1635444444
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1635444444
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_97
timestamp 1635444444
transform 1 0 10028 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1635444444
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_7
timestamp 1635444444
transform 1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1635444444
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1635444444
transform -1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1635444444
transform -1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_15
timestamp 1635444444
transform 1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_22
timestamp 1635444444
transform 1 0 3128 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _109_
timestamp 1635444444
transform 1 0 2852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_29
timestamp 1635444444
transform 1 0 3772 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1635444444
transform -1 0 3772 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_41
timestamp 1635444444
transform 1 0 4876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1635444444
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1635444444
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1635444444
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1635444444
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_93
timestamp 1635444444
transform 1 0 9660 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_99
timestamp 1635444444
transform 1 0 10212 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1635444444
transform 1 0 9844 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1635444444
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_84_7
timestamp 1635444444
transform 1 0 1748 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1635444444
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1635444444
transform -1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_15
timestamp 1635444444
transform 1 0 2484 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_19
timestamp 1635444444
transform 1 0 2852 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _216_
timestamp 1635444444
transform -1 0 2852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1635444444
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1635444444
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1635444444
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1635444444
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1635444444
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1635444444
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1635444444
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_85
timestamp 1635444444
transform 1 0 8924 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_93
timestamp 1635444444
transform 1 0 9660 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_99
timestamp 1635444444
transform 1 0 10212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1635444444
transform 1 0 9844 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1635444444
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_7
timestamp 1635444444
transform 1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_10
timestamp 1635444444
transform 1 0 2024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1635444444
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1635444444
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1635444444
transform -1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1635444444
transform -1 0 2484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1635444444
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_18
timestamp 1635444444
transform 1 0 2760 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1635444444
transform 1 0 2392 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1635444444
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_26
timestamp 1635444444
transform 1 0 3496 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_35
timestamp 1635444444
transform 1 0 4324 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  _200_
timestamp 1635444444
transform 1 0 3772 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1635444444
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1635444444
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_47
timestamp 1635444444
transform 1 0 5428 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1635444444
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1635444444
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_59
timestamp 1635444444
transform 1 0 6532 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1635444444
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_71
timestamp 1635444444
transform 1 0 7636 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1635444444
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1635444444
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_85
timestamp 1635444444
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_101
timestamp 1635444444
transform 1 0 10396 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_85_93
timestamp 1635444444
transform 1 0 9660 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_93
timestamp 1635444444
transform 1 0 9660 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_99
timestamp 1635444444
transform 1 0 10212 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1635444444
transform 1 0 9844 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1635444444
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1635444444
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_10
timestamp 1635444444
transform 1 0 2024 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1635444444
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _146_
timestamp 1635444444
transform -1 0 2024 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_87_18
timestamp 1635444444
transform 1 0 2760 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1635444444
transform 1 0 2392 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_30
timestamp 1635444444
transform 1 0 3864 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_42
timestamp 1635444444
transform 1 0 4968 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_54
timestamp 1635444444
transform 1 0 6072 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1635444444
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1635444444
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1635444444
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_93
timestamp 1635444444
transform 1 0 9660 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_99
timestamp 1635444444
transform 1 0 10212 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1635444444
transform 1 0 9844 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1635444444
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1635444444
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1635444444
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _147_
timestamp 1635444444
transform -1 0 2024 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_88_17
timestamp 1635444444
transform 1 0 2668 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_24
timestamp 1635444444
transform 1 0 3312 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _125_
timestamp 1635444444
transform -1 0 2668 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _127_
timestamp 1635444444
transform 1 0 3036 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_32
timestamp 1635444444
transform 1 0 4048 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 1635444444
transform -1 0 4048 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_44
timestamp 1635444444
transform 1 0 5152 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_56
timestamp 1635444444
transform 1 0 6256 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_68
timestamp 1635444444
transform 1 0 7360 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_80
timestamp 1635444444
transform 1 0 8464 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_88_85
timestamp 1635444444
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_93
timestamp 1635444444
transform 1 0 9660 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_99
timestamp 1635444444
transform 1 0 10212 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1635444444
transform 1 0 9844 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1635444444
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_7
timestamp 1635444444
transform 1 0 1748 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1635444444
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1635444444
transform -1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_19
timestamp 1635444444
transform 1 0 2852 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_24
timestamp 1635444444
transform 1 0 3312 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _218_
timestamp 1635444444
transform 1 0 3036 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_36
timestamp 1635444444
transform 1 0 4416 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_48
timestamp 1635444444
transform 1 0 5520 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1635444444
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1635444444
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1635444444
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_101
timestamp 1635444444
transform 1 0 10396 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_93
timestamp 1635444444
transform 1 0 9660 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1635444444
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_7
timestamp 1635444444
transform 1 0 1748 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1635444444
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1635444444
transform -1 0 1748 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1635444444
transform -1 0 2484 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_15
timestamp 1635444444
transform 1 0 2484 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_23
timestamp 1635444444
transform 1 0 3220 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1635444444
transform 1 0 2852 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1635444444
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1635444444
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1635444444
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1635444444
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1635444444
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1635444444
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1635444444
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_85
timestamp 1635444444
transform 1 0 8924 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_93
timestamp 1635444444
transform 1 0 9660 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_99
timestamp 1635444444
transform 1 0 10212 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1635444444
transform 1 0 9844 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1635444444
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_10
timestamp 1635444444
transform 1 0 2024 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1635444444
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _144_
timestamp 1635444444
transform 1 0 1380 0 -1 52224
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_91_17
timestamp 1635444444
transform 1 0 2668 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_91_24
timestamp 1635444444
transform 1 0 3312 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _129_
timestamp 1635444444
transform -1 0 2668 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _219_
timestamp 1635444444
transform -1 0 3312 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_36
timestamp 1635444444
transform 1 0 4416 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_48
timestamp 1635444444
transform 1 0 5520 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1635444444
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1635444444
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1635444444
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_93
timestamp 1635444444
transform 1 0 9660 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_99
timestamp 1635444444
transform 1 0 10212 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1635444444
transform 1 0 9844 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1635444444
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_92_11
timestamp 1635444444
transform 1 0 2116 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_7
timestamp 1635444444
transform 1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_7
timestamp 1635444444
transform 1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1635444444
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1635444444
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _111_
timestamp 1635444444
transform 1 0 2208 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1635444444
transform -1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1635444444
transform -1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1635444444
transform 1 0 2116 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1635444444
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_15
timestamp 1635444444
transform 1 0 2484 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_23
timestamp 1635444444
transform 1 0 3220 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1635444444
transform 1 0 2852 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1635444444
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1635444444
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_35
timestamp 1635444444
transform 1 0 4324 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1635444444
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1635444444
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1635444444
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1635444444
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1635444444
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1635444444
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1635444444
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1635444444
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1635444444
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_85
timestamp 1635444444
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1635444444
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_97
timestamp 1635444444
transform 1 0 10028 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_93
timestamp 1635444444
transform 1 0 9660 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_99
timestamp 1635444444
transform 1 0 10212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1635444444
transform 1 0 9844 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1635444444
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1635444444
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_11
timestamp 1635444444
transform 1 0 2116 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1635444444
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _143_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_94_18
timestamp 1635444444
transform 1 0 2760 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _131_
timestamp 1635444444
transform -1 0 2760 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1635444444
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1635444444
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1635444444
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1635444444
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1635444444
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1635444444
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1635444444
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_85
timestamp 1635444444
transform 1 0 8924 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_93
timestamp 1635444444
transform 1 0 9660 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_99
timestamp 1635444444
transform 1 0 10212 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1635444444
transform 1 0 9844 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1635444444
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_7
timestamp 1635444444
transform 1 0 1748 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1635444444
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1635444444
transform -1 0 1748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_15
timestamp 1635444444
transform 1 0 2484 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_21
timestamp 1635444444
transform 1 0 3036 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _220_
timestamp 1635444444
transform -1 0 3036 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_33
timestamp 1635444444
transform 1 0 4140 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_45
timestamp 1635444444
transform 1 0 5244 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_53
timestamp 1635444444
transform 1 0 5980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1635444444
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1635444444
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1635444444
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_93
timestamp 1635444444
transform 1 0 9660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1635444444
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1635444444
transform 1 0 9844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1635444444
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_7
timestamp 1635444444
transform 1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1635444444
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1635444444
transform -1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1635444444
transform 1 0 2116 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1635444444
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1635444444
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1635444444
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1635444444
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1635444444
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1635444444
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1635444444
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1635444444
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_85
timestamp 1635444444
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_97
timestamp 1635444444
transform 1 0 10028 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1635444444
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_97_10
timestamp 1635444444
transform 1 0 2024 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1635444444
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _149_
timestamp 1635444444
transform 1 0 1380 0 -1 55488
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_8  _104_
timestamp 1635444444
transform 1 0 2576 0 -1 55488
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1635444444
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1635444444
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1635444444
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1635444444
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1635444444
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1635444444
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1635444444
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_93
timestamp 1635444444
transform 1 0 9660 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_99
timestamp 1635444444
transform 1 0 10212 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635444444
transform 1 0 9936 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1635444444
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_7
timestamp 1635444444
transform 1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1635444444
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1635444444
transform -1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1635444444
transform 1 0 2116 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_15
timestamp 1635444444
transform 1 0 2484 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_22
timestamp 1635444444
transform 1 0 3128 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1635444444
transform -1 0 3128 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_29
timestamp 1635444444
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_41
timestamp 1635444444
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_53
timestamp 1635444444
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_65
timestamp 1635444444
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1635444444
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1635444444
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_85
timestamp 1635444444
transform 1 0 8924 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_98_93
timestamp 1635444444
transform 1 0 9660 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_99
timestamp 1635444444
transform 1 0 10212 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635444444
transform 1 0 9936 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1635444444
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_100_7
timestamp 1635444444
transform 1 0 1748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_7
timestamp 1635444444
transform 1 0 1748 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1635444444
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1635444444
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1635444444
transform -1 0 1748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1635444444
transform -1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1635444444
transform -1 0 2484 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_15
timestamp 1635444444
transform 1 0 2484 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_22
timestamp 1635444444
transform 1 0 3128 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_13
timestamp 1635444444
transform 1 0 2300 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_20
timestamp 1635444444
transform 1 0 2944 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _133_
timestamp 1635444444
transform -1 0 3128 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _141_
timestamp 1635444444
transform -1 0 2944 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _222_
timestamp 1635444444
transform -1 0 3588 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_32
timestamp 1635444444
transform 1 0 4048 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1635444444
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _221_
timestamp 1635444444
transform -1 0 4048 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_44
timestamp 1635444444
transform 1 0 5152 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1635444444
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1635444444
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_56
timestamp 1635444444
transform 1 0 6256 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1635444444
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1635444444
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_68
timestamp 1635444444
transform 1 0 7360 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1635444444
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_80
timestamp 1635444444
transform 1 0 8464 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_85
timestamp 1635444444
transform 1 0 8924 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1635444444
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1635444444
transform -1 0 10212 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1635444444
transform 1 0 10212 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_101
timestamp 1635444444
transform 1 0 10396 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_93
timestamp 1635444444
transform 1 0 9660 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1635444444
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1635444444
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_7
timestamp 1635444444
transform 1 0 1748 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1635444444
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1635444444
transform -1 0 1748 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1635444444
transform -1 0 2484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_15
timestamp 1635444444
transform 1 0 2484 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_101_22
timestamp 1635444444
transform 1 0 3128 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _135_
timestamp 1635444444
transform 1 0 2852 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_34
timestamp 1635444444
transform 1 0 4232 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_46
timestamp 1635444444
transform 1 0 5336 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1635444444
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1635444444
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1635444444
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_81
timestamp 1635444444
transform 1 0 8556 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1635444444
transform -1 0 10212 0 -1 57664
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_101_99
timestamp 1635444444
transform 1 0 10212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1635444444
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_12
timestamp 1635444444
transform 1 0 2208 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_3
timestamp 1635444444
transform 1 0 1380 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1635444444
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _148_
timestamp 1635444444
transform 1 0 1472 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_102_20
timestamp 1635444444
transform 1 0 2944 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1635444444
transform 1 0 2576 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_32
timestamp 1635444444
transform 1 0 4048 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1635444444
transform -1 0 4048 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_102_44
timestamp 1635444444
transform 1 0 5152 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_56
timestamp 1635444444
transform 1 0 6256 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_68
timestamp 1635444444
transform 1 0 7360 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_102_80
timestamp 1635444444
transform 1 0 8464 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_102_85
timestamp 1635444444
transform 1 0 8924 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_102_97
timestamp 1635444444
transform 1 0 10028 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1635444444
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_103_12
timestamp 1635444444
transform 1 0 2208 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_3
timestamp 1635444444
transform 1 0 1380 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1635444444
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _153_
timestamp 1635444444
transform -1 0 2208 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_103_20
timestamp 1635444444
transform 1 0 2944 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1635444444
transform 1 0 2576 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_32
timestamp 1635444444
transform 1 0 4048 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_44
timestamp 1635444444
transform 1 0 5152 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1635444444
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1635444444
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_81
timestamp 1635444444
transform 1 0 8556 0 -1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1635444444
transform -1 0 10212 0 -1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1635444444
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1635444444
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_11
timestamp 1635444444
transform 1 0 2116 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1635444444
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _150_
timestamp 1635444444
transform 1 0 1380 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_104_19
timestamp 1635444444
transform 1 0 2852 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1635444444
transform -1 0 2852 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1635444444
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1635444444
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1635444444
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1635444444
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1635444444
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1635444444
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1635444444
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_85
timestamp 1635444444
transform 1 0 8924 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_93
timestamp 1635444444
transform 1 0 9660 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_99
timestamp 1635444444
transform 1 0 10212 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 9936 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1635444444
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_7
timestamp 1635444444
transform 1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_3
timestamp 1635444444
transform 1 0 1380 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_9
timestamp 1635444444
transform 1 0 1932 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1635444444
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1635444444
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _151_
timestamp 1635444444
transform 1 0 2024 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _152_
timestamp 1635444444
transform 1 0 2116 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1635444444
transform -1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_19
timestamp 1635444444
transform 1 0 2852 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_106_18
timestamp 1635444444
transform 1 0 2760 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1635444444
transform 1 0 3220 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1635444444
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_26
timestamp 1635444444
transform 1 0 3496 0 1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1635444444
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1635444444
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1635444444
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1635444444
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1635444444
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1635444444
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1635444444
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1635444444
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1635444444
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1635444444
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1635444444
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1635444444
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_85
timestamp 1635444444
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_105_93
timestamp 1635444444
transform 1 0 9660 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_99
timestamp 1635444444
transform 1 0 10212 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_97
timestamp 1635444444
transform 1 0 10028 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 9936 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1635444444
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1635444444
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_12
timestamp 1635444444
transform 1 0 2208 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_3
timestamp 1635444444
transform 1 0 1380 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1635444444
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _154_
timestamp 1635444444
transform 1 0 1472 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_20
timestamp 1635444444
transform 1 0 2944 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1635444444
transform 1 0 2576 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_32
timestamp 1635444444
transform 1 0 4048 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_44
timestamp 1635444444
transform 1 0 5152 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1635444444
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1635444444
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1635444444
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_93
timestamp 1635444444
transform 1 0 9660 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1635444444
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635444444
transform 1 0 9936 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1635444444
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_108_7
timestamp 1635444444
transform 1 0 1748 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1635444444
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1635444444
transform -1 0 1748 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_13
timestamp 1635444444
transform 1 0 2300 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_21
timestamp 1635444444
transform 1 0 3036 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _176_
timestamp 1635444444
transform 1 0 2392 0 1 60928
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1635444444
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_29
timestamp 1635444444
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_41
timestamp 1635444444
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_53
timestamp 1635444444
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_65
timestamp 1635444444
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1635444444
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1635444444
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_85
timestamp 1635444444
transform 1 0 8924 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_108_93
timestamp 1635444444
transform 1 0 9660 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_99
timestamp 1635444444
transform 1 0 10212 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635444444
transform 1 0 9936 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1635444444
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_7
timestamp 1635444444
transform 1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1635444444
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1635444444
transform -1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1635444444
transform -1 0 2484 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1635444444
transform 1 0 2484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1635444444
transform 1 0 3588 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_39
timestamp 1635444444
transform 1 0 4692 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_51
timestamp 1635444444
transform 1 0 5796 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1635444444
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1635444444
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1635444444
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1635444444
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_109_101
timestamp 1635444444
transform 1 0 10396 0 -1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_109_93
timestamp 1635444444
transform 1 0 9660 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1635444444
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_110_7
timestamp 1635444444
transform 1 0 1748 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1635444444
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1635444444
transform -1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_110_21
timestamp 1635444444
transform 1 0 3036 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _159_
timestamp 1635444444
transform -1 0 3036 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1635444444
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1635444444
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1635444444
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1635444444
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1635444444
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1635444444
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1635444444
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_85
timestamp 1635444444
transform 1 0 8924 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_110_93
timestamp 1635444444
transform 1 0 9660 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_99
timestamp 1635444444
transform 1 0 10212 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635444444
transform 1 0 9936 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1635444444
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_111_11
timestamp 1635444444
transform 1 0 2116 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1635444444
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _155_
timestamp 1635444444
transform 1 0 1380 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_23
timestamp 1635444444
transform 1 0 3220 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _139_
timestamp 1635444444
transform -1 0 3220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_111_35
timestamp 1635444444
transform 1 0 4324 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_111_47
timestamp 1635444444
transform 1 0 5428 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1635444444
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1635444444
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1635444444
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1635444444
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_93
timestamp 1635444444
transform 1 0 9660 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_99
timestamp 1635444444
transform 1 0 10212 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635444444
transform 1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1635444444
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_7
timestamp 1635444444
transform 1 0 1748 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_7
timestamp 1635444444
transform 1 0 1748 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1635444444
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1635444444
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1635444444
transform -1 0 1748 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1635444444
transform -1 0 1748 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1635444444
transform 1 0 2116 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1635444444
transform -1 0 2484 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_15
timestamp 1635444444
transform 1 0 2484 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_112_23
timestamp 1635444444
transform 1 0 3220 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1635444444
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1635444444
transform 1 0 2852 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1635444444
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_29
timestamp 1635444444
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1635444444
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_41
timestamp 1635444444
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_39
timestamp 1635444444
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1635444444
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_53
timestamp 1635444444
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1635444444
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1635444444
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_65
timestamp 1635444444
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1635444444
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1635444444
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1635444444
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_85
timestamp 1635444444
transform 1 0 8924 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_113_81
timestamp 1635444444
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_112_93
timestamp 1635444444
transform 1 0 9660 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_99
timestamp 1635444444
transform 1 0 10212 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_113_101
timestamp 1635444444
transform 1 0 10396 0 -1 64192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_113_93
timestamp 1635444444
transform 1 0 9660 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635444444
transform 1 0 9936 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1635444444
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1635444444
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_11
timestamp 1635444444
transform 1 0 2116 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1635444444
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _156_
timestamp 1635444444
transform 1 0 1380 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_114_19
timestamp 1635444444
transform 1 0 2852 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1635444444
transform 1 0 2484 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1635444444
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1635444444
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1635444444
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1635444444
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1635444444
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1635444444
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1635444444
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_85
timestamp 1635444444
transform 1 0 8924 0 1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_114_93
timestamp 1635444444
transform 1 0 9660 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_114_99
timestamp 1635444444
transform 1 0 10212 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1635444444
transform 1 0 9936 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1635444444
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_115_10
timestamp 1635444444
transform 1 0 2024 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1635444444
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _142_
timestamp 1635444444
transform 1 0 1380 0 -1 65280
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_115_24
timestamp 1635444444
transform 1 0 3312 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _158_
timestamp 1635444444
transform -1 0 3312 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_115_32
timestamp 1635444444
transform 1 0 4048 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1635444444
transform 1 0 3680 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_115_44
timestamp 1635444444
transform 1 0 5152 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1635444444
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1635444444
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1635444444
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_93
timestamp 1635444444
transform 1 0 9660 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_99
timestamp 1635444444
transform 1 0 10212 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1635444444
transform 1 0 9936 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1635444444
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_6
timestamp 1635444444
transform 1 0 1656 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1635444444
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _160_
timestamp 1635444444
transform -1 0 2760 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1635444444
transform -1 0 1656 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_116_18
timestamp 1635444444
transform 1 0 2760 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_116_26
timestamp 1635444444
transform 1 0 3496 0 1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_116_33
timestamp 1635444444
transform 1 0 4140 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1635444444
transform 1 0 3772 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_45
timestamp 1635444444
transform 1 0 5244 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_57
timestamp 1635444444
transform 1 0 6348 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_69
timestamp 1635444444
transform 1 0 7452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_116_81
timestamp 1635444444
transform 1 0 8556 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_116_85
timestamp 1635444444
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_116_97
timestamp 1635444444
transform 1 0 10028 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1635444444
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_11
timestamp 1635444444
transform 1 0 2116 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1635444444
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _157_
timestamp 1635444444
transform 1 0 1380 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_23
timestamp 1635444444
transform 1 0 3220 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _161_
timestamp 1635444444
transform 1 0 2484 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_117_35
timestamp 1635444444
transform 1 0 4324 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_47
timestamp 1635444444
transform 1 0 5428 0 -1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1635444444
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1635444444
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1635444444
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1635444444
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_93
timestamp 1635444444
transform 1 0 9660 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1635444444
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635444444
transform 1 0 9936 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1635444444
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1635444444
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1635444444
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1635444444
transform 1 0 1380 0 1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1635444444
transform 1 0 1380 0 -1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_118_13
timestamp 1635444444
transform 1 0 2300 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_118_21
timestamp 1635444444
transform 1 0 3036 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_13
timestamp 1635444444
transform 1 0 2300 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_25
timestamp 1635444444
transform 1 0 3404 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1635444444
transform -1 0 3036 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1635444444
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1635444444
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_37
timestamp 1635444444
transform 1 0 4508 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1635444444
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_49
timestamp 1635444444
transform 1 0 5612 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1635444444
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1635444444
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1635444444
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1635444444
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1635444444
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1635444444
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1635444444
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_85
timestamp 1635444444
transform 1 0 8924 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1635444444
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_118_93
timestamp 1635444444
transform 1 0 9660 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_99
timestamp 1635444444
transform 1 0 10212 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_119_93
timestamp 1635444444
transform 1 0 9660 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_119_99
timestamp 1635444444
transform 1 0 10212 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635444444
transform 1 0 9936 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635444444
transform 1 0 9936 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1635444444
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1635444444
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1635444444
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1635444444
transform 1 0 1380 0 1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_120_13
timestamp 1635444444
transform 1 0 2300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_120_25
timestamp 1635444444
transform 1 0 3404 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1635444444
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1635444444
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1635444444
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1635444444
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1635444444
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1635444444
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_85
timestamp 1635444444
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_120_97
timestamp 1635444444
transform 1 0 10028 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1635444444
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1635444444
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1635444444
transform 1 0 1380 0 -1 68544
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_121_13
timestamp 1635444444
transform 1 0 2300 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_25
timestamp 1635444444
transform 1 0 3404 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _162_
timestamp 1635444444
transform 1 0 2668 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_121_37
timestamp 1635444444
transform 1 0 4508 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_49
timestamp 1635444444
transform 1 0 5612 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1635444444
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1635444444
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1635444444
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1635444444
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_93
timestamp 1635444444
transform 1 0 9660 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_99
timestamp 1635444444
transform 1 0 10212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635444444
transform 1 0 9936 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1635444444
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_122_6
timestamp 1635444444
transform 1 0 1656 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1635444444
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _168_
timestamp 1635444444
transform -1 0 2944 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635444444
transform -1 0 1656 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_20
timestamp 1635444444
transform 1 0 2944 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_29
timestamp 1635444444
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_41
timestamp 1635444444
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_53
timestamp 1635444444
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_65
timestamp 1635444444
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1635444444
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1635444444
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_85
timestamp 1635444444
transform 1 0 8924 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_122_93
timestamp 1635444444
transform 1 0 9660 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_99
timestamp 1635444444
transform 1 0 10212 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635444444
transform 1 0 9936 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1635444444
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_123_11
timestamp 1635444444
transform 1 0 2116 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1635444444
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _163_
timestamp 1635444444
transform 1 0 1380 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_123_18
timestamp 1635444444
transform 1 0 2760 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_25
timestamp 1635444444
transform 1 0 3404 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635444444
transform 1 0 2484 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635444444
transform 1 0 3128 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_37
timestamp 1635444444
transform 1 0 4508 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_49
timestamp 1635444444
transform 1 0 5612 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1635444444
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1635444444
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1635444444
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1635444444
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_123_101
timestamp 1635444444
transform 1 0 10396 0 -1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_123_93
timestamp 1635444444
transform 1 0 9660 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1635444444
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_11
timestamp 1635444444
transform 1 0 2116 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1635444444
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _164_
timestamp 1635444444
transform 1 0 1380 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_124_18
timestamp 1635444444
transform 1 0 2760 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform 1 0 2484 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_124_26
timestamp 1635444444
transform 1 0 3496 0 1 69632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_124_29
timestamp 1635444444
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_41
timestamp 1635444444
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_53
timestamp 1635444444
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_65
timestamp 1635444444
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1635444444
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1635444444
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_85
timestamp 1635444444
transform 1 0 8924 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_124_93
timestamp 1635444444
transform 1 0 9660 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1635444444
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform 1 0 9936 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1635444444
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_11
timestamp 1635444444
transform 1 0 2116 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_6
timestamp 1635444444
transform 1 0 1656 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1635444444
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1635444444
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _165_
timestamp 1635444444
transform 1 0 1380 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _169_
timestamp 1635444444
transform 1 0 2208 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform -1 0 1656 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_18
timestamp 1635444444
transform 1 0 2760 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_20
timestamp 1635444444
transform 1 0 2944 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform 1 0 2484 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_30
timestamp 1635444444
transform 1 0 3864 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1635444444
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_42
timestamp 1635444444
transform 1 0 4968 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1635444444
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_125_54
timestamp 1635444444
transform 1 0 6072 0 -1 70720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1635444444
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1635444444
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1635444444
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1635444444
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1635444444
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1635444444
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1635444444
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1635444444
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_125_93
timestamp 1635444444
transform 1 0 9660 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_99
timestamp 1635444444
transform 1 0 10212 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_97
timestamp 1635444444
transform 1 0 10028 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635444444
transform 1 0 9936 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1635444444
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1635444444
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_6
timestamp 1635444444
transform 1 0 1656 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1635444444
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1635444444
transform -1 0 1656 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1635444444
transform 1 0 2024 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_13
timestamp 1635444444
transform 1 0 2300 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_25
timestamp 1635444444
transform 1 0 3404 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_37
timestamp 1635444444
transform 1 0 4508 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_49
timestamp 1635444444
transform 1 0 5612 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1635444444
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1635444444
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1635444444
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1635444444
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_93
timestamp 1635444444
transform 1 0 9660 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_99
timestamp 1635444444
transform 1 0 10212 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635444444
transform 1 0 9936 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1635444444
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_6
timestamp 1635444444
transform 1 0 1656 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1635444444
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1635444444
transform -1 0 1656 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform -1 0 2300 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_13
timestamp 1635444444
transform 1 0 2300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_128_25
timestamp 1635444444
transform 1 0 3404 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1635444444
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1635444444
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1635444444
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1635444444
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1635444444
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1635444444
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_85
timestamp 1635444444
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_128_93
timestamp 1635444444
transform 1 0 9660 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1635444444
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635444444
transform 1 0 9936 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1635444444
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_129_6
timestamp 1635444444
transform 1 0 1656 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1635444444
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _170_
timestamp 1635444444
transform -1 0 2944 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform -1 0 1656 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_20
timestamp 1635444444
transform 1 0 2944 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_32
timestamp 1635444444
transform 1 0 4048 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_44
timestamp 1635444444
transform 1 0 5152 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1635444444
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1635444444
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1635444444
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_129_93
timestamp 1635444444
transform 1 0 9660 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_129_99
timestamp 1635444444
transform 1 0 10212 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1635444444
transform 1 0 9936 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1635444444
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_11
timestamp 1635444444
transform 1 0 2116 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1635444444
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _167_
timestamp 1635444444
transform -1 0 2116 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_130_18
timestamp 1635444444
transform 1 0 2760 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform -1 0 2760 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_130_26
timestamp 1635444444
transform 1 0 3496 0 1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1635444444
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1635444444
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1635444444
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1635444444
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1635444444
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1635444444
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_85
timestamp 1635444444
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_130_97
timestamp 1635444444
transform 1 0 10028 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1635444444
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_11
timestamp 1635444444
transform 1 0 2116 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1635444444
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _166_
timestamp 1635444444
transform -1 0 2116 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_18
timestamp 1635444444
transform 1 0 2760 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635444444
transform 1 0 2484 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_30
timestamp 1635444444
transform 1 0 3864 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_42
timestamp 1635444444
transform 1 0 4968 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_54
timestamp 1635444444
transform 1 0 6072 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1635444444
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1635444444
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1635444444
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_93
timestamp 1635444444
transform 1 0 9660 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_99
timestamp 1635444444
transform 1 0 10212 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635444444
transform 1 0 9936 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1635444444
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_6
timestamp 1635444444
transform 1 0 1656 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_6
timestamp 1635444444
transform 1 0 1656 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1635444444
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1635444444
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _171_
timestamp 1635444444
transform -1 0 2944 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform -1 0 1656 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1635444444
transform -1 0 1656 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_132_18
timestamp 1635444444
transform 1 0 2760 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_20
timestamp 1635444444
transform 1 0 2944 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_132_26
timestamp 1635444444
transform 1 0 3496 0 1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1635444444
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_32
timestamp 1635444444
transform 1 0 4048 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1635444444
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_44
timestamp 1635444444
transform 1 0 5152 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_53
timestamp 1635444444
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1635444444
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_65
timestamp 1635444444
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1635444444
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1635444444
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1635444444
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_85
timestamp 1635444444
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1635444444
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_132_93
timestamp 1635444444
transform 1 0 9660 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1635444444
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_133_101
timestamp 1635444444
transform 1 0 10396 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_133_93
timestamp 1635444444
transform 1 0 9660 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635444444
transform 1 0 9936 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1635444444
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1635444444
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_3
timestamp 1635444444
transform 1 0 1380 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_134_7
timestamp 1635444444
transform 1 0 1748 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1635444444
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _173_
timestamp 1635444444
transform 1 0 1840 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_134_16
timestamp 1635444444
transform 1 0 2576 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_134_23
timestamp 1635444444
transform 1 0 3220 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform 1 0 2944 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1635444444
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_29
timestamp 1635444444
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_41
timestamp 1635444444
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_53
timestamp 1635444444
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_65
timestamp 1635444444
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1635444444
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1635444444
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1635444444
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_134_93
timestamp 1635444444
transform 1 0 9660 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1635444444
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635444444
transform 1 0 9936 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1635444444
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_135_12
timestamp 1635444444
transform 1 0 2208 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_135_6
timestamp 1635444444
transform 1 0 1656 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1635444444
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform -1 0 1656 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_21
timestamp 1635444444
transform 1 0 3036 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _172_
timestamp 1635444444
transform 1 0 2300 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform 1 0 3404 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_28
timestamp 1635444444
transform 1 0 3680 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_40
timestamp 1635444444
transform 1 0 4784 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_52
timestamp 1635444444
transform 1 0 5888 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1635444444
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1635444444
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1635444444
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_135_93
timestamp 1635444444
transform 1 0 9660 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_99
timestamp 1635444444
transform 1 0 10212 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635444444
transform 1 0 9936 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1635444444
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_3
timestamp 1635444444
transform 1 0 1380 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_7
timestamp 1635444444
transform 1 0 1748 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1635444444
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _174_
timestamp 1635444444
transform 1 0 1840 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_136_16
timestamp 1635444444
transform 1 0 2576 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_136_23
timestamp 1635444444
transform 1 0 3220 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform 1 0 2944 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1635444444
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_32
timestamp 1635444444
transform 1 0 4048 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1635444444
transform 1 0 3772 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_44
timestamp 1635444444
transform 1 0 5152 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_56
timestamp 1635444444
transform 1 0 6256 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_68
timestamp 1635444444
transform 1 0 7360 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_80
timestamp 1635444444
transform 1 0 8464 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_136_85
timestamp 1635444444
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_136_93
timestamp 1635444444
transform 1 0 9660 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1635444444
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1635444444
transform 1 0 9936 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1635444444
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_11
timestamp 1635444444
transform 1 0 2116 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1635444444
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _175_
timestamp 1635444444
transform 1 0 1380 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_137_18
timestamp 1635444444
transform 1 0 2760 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_25
timestamp 1635444444
transform 1 0 3404 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform 1 0 2484 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform 1 0 3128 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_32
timestamp 1635444444
transform 1 0 4048 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform 1 0 3772 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform 1 0 4416 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_39
timestamp 1635444444
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1635444444
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1635444444
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1635444444
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1635444444
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_81
timestamp 1635444444
transform 1 0 8556 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_87
timestamp 1635444444
transform 1 0 9108 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1635444444
transform 1 0 9200 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_91
timestamp 1635444444
transform 1 0 9476 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1635444444
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1635444444
transform -1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1635444444
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1635444444
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1635444444
transform 1 0 1380 0 1 77248
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_138_13
timestamp 1635444444
transform 1 0 2300 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_20
timestamp 1635444444
transform 1 0 2944 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1635444444
transform 1 0 2668 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_32
timestamp 1635444444
transform 1 0 4048 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform 1 0 3772 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform 1 0 4416 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_39
timestamp 1635444444
transform 1 0 4692 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_51
timestamp 1635444444
transform 1 0 5796 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_138_55
timestamp 1635444444
transform 1 0 6164 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1635444444
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1635444444
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1635444444
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_138_85
timestamp 1635444444
transform 1 0 8924 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635444444
transform 1 0 9200 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_91
timestamp 1635444444
transform 1 0 9476 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1635444444
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1635444444
transform -1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1635444444
transform -1 0 10856 0 1 77248
box -38 -48 314 592
<< labels >>
rlabel metal4 s 2575 2128 2895 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 5839 2128 6159 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 9103 2128 9423 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 4207 2128 4527 77840 6 vssd1
port 1 nsew ground input
rlabel metal4 s 7471 2128 7791 77840 6 vssd1
port 1 nsew ground input
rlabel metal2 s 2962 0 3018 800 6 wb_clk_i
port 2 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wb_rst_i
port 3 nsew signal input
rlabel metal3 s 11200 79432 12000 79552 6 wbm_a_ack_i
port 4 nsew signal input
rlabel metal3 s 11200 5584 12000 5704 6 wbm_a_adr_o[0]
port 5 nsew signal tristate
rlabel metal3 s 11200 13336 12000 13456 6 wbm_a_adr_o[10]
port 6 nsew signal tristate
rlabel metal3 s 11200 14016 12000 14136 6 wbm_a_adr_o[11]
port 7 nsew signal tristate
rlabel metal3 s 11200 14832 12000 14952 6 wbm_a_adr_o[12]
port 8 nsew signal tristate
rlabel metal3 s 11200 15648 12000 15768 6 wbm_a_adr_o[13]
port 9 nsew signal tristate
rlabel metal3 s 11200 16328 12000 16448 6 wbm_a_adr_o[14]
port 10 nsew signal tristate
rlabel metal3 s 11200 17144 12000 17264 6 wbm_a_adr_o[15]
port 11 nsew signal tristate
rlabel metal3 s 11200 17960 12000 18080 6 wbm_a_adr_o[16]
port 12 nsew signal tristate
rlabel metal3 s 11200 18640 12000 18760 6 wbm_a_adr_o[17]
port 13 nsew signal tristate
rlabel metal3 s 11200 19456 12000 19576 6 wbm_a_adr_o[18]
port 14 nsew signal tristate
rlabel metal3 s 11200 20272 12000 20392 6 wbm_a_adr_o[19]
port 15 nsew signal tristate
rlabel metal3 s 11200 6400 12000 6520 6 wbm_a_adr_o[1]
port 16 nsew signal tristate
rlabel metal3 s 11200 20952 12000 21072 6 wbm_a_adr_o[20]
port 17 nsew signal tristate
rlabel metal3 s 11200 21768 12000 21888 6 wbm_a_adr_o[21]
port 18 nsew signal tristate
rlabel metal3 s 11200 22448 12000 22568 6 wbm_a_adr_o[22]
port 19 nsew signal tristate
rlabel metal3 s 11200 23264 12000 23384 6 wbm_a_adr_o[23]
port 20 nsew signal tristate
rlabel metal3 s 11200 24080 12000 24200 6 wbm_a_adr_o[24]
port 21 nsew signal tristate
rlabel metal3 s 11200 24760 12000 24880 6 wbm_a_adr_o[25]
port 22 nsew signal tristate
rlabel metal3 s 11200 25576 12000 25696 6 wbm_a_adr_o[26]
port 23 nsew signal tristate
rlabel metal3 s 11200 26392 12000 26512 6 wbm_a_adr_o[27]
port 24 nsew signal tristate
rlabel metal3 s 11200 27072 12000 27192 6 wbm_a_adr_o[28]
port 25 nsew signal tristate
rlabel metal3 s 11200 27888 12000 28008 6 wbm_a_adr_o[29]
port 26 nsew signal tristate
rlabel metal3 s 11200 7080 12000 7200 6 wbm_a_adr_o[2]
port 27 nsew signal tristate
rlabel metal3 s 11200 28704 12000 28824 6 wbm_a_adr_o[30]
port 28 nsew signal tristate
rlabel metal3 s 11200 29384 12000 29504 6 wbm_a_adr_o[31]
port 29 nsew signal tristate
rlabel metal3 s 11200 7896 12000 8016 6 wbm_a_adr_o[3]
port 30 nsew signal tristate
rlabel metal3 s 11200 8712 12000 8832 6 wbm_a_adr_o[4]
port 31 nsew signal tristate
rlabel metal3 s 11200 9392 12000 9512 6 wbm_a_adr_o[5]
port 32 nsew signal tristate
rlabel metal3 s 11200 10208 12000 10328 6 wbm_a_adr_o[6]
port 33 nsew signal tristate
rlabel metal3 s 11200 11024 12000 11144 6 wbm_a_adr_o[7]
port 34 nsew signal tristate
rlabel metal3 s 11200 11704 12000 11824 6 wbm_a_adr_o[8]
port 35 nsew signal tristate
rlabel metal3 s 11200 12520 12000 12640 6 wbm_a_adr_o[9]
port 36 nsew signal tristate
rlabel metal3 s 11200 960 12000 1080 6 wbm_a_cyc_o
port 37 nsew signal tristate
rlabel metal3 s 11200 54816 12000 54936 6 wbm_a_dat_i[0]
port 38 nsew signal input
rlabel metal3 s 11200 62432 12000 62552 6 wbm_a_dat_i[10]
port 39 nsew signal input
rlabel metal3 s 11200 63248 12000 63368 6 wbm_a_dat_i[11]
port 40 nsew signal input
rlabel metal3 s 11200 64064 12000 64184 6 wbm_a_dat_i[12]
port 41 nsew signal input
rlabel metal3 s 11200 64744 12000 64864 6 wbm_a_dat_i[13]
port 42 nsew signal input
rlabel metal3 s 11200 65560 12000 65680 6 wbm_a_dat_i[14]
port 43 nsew signal input
rlabel metal3 s 11200 66376 12000 66496 6 wbm_a_dat_i[15]
port 44 nsew signal input
rlabel metal3 s 11200 67056 12000 67176 6 wbm_a_dat_i[16]
port 45 nsew signal input
rlabel metal3 s 11200 67872 12000 67992 6 wbm_a_dat_i[17]
port 46 nsew signal input
rlabel metal3 s 11200 68688 12000 68808 6 wbm_a_dat_i[18]
port 47 nsew signal input
rlabel metal3 s 11200 69368 12000 69488 6 wbm_a_dat_i[19]
port 48 nsew signal input
rlabel metal3 s 11200 55632 12000 55752 6 wbm_a_dat_i[1]
port 49 nsew signal input
rlabel metal3 s 11200 70184 12000 70304 6 wbm_a_dat_i[20]
port 50 nsew signal input
rlabel metal3 s 11200 71000 12000 71120 6 wbm_a_dat_i[21]
port 51 nsew signal input
rlabel metal3 s 11200 71680 12000 71800 6 wbm_a_dat_i[22]
port 52 nsew signal input
rlabel metal3 s 11200 72496 12000 72616 6 wbm_a_dat_i[23]
port 53 nsew signal input
rlabel metal3 s 11200 73312 12000 73432 6 wbm_a_dat_i[24]
port 54 nsew signal input
rlabel metal3 s 11200 73992 12000 74112 6 wbm_a_dat_i[25]
port 55 nsew signal input
rlabel metal3 s 11200 74808 12000 74928 6 wbm_a_dat_i[26]
port 56 nsew signal input
rlabel metal3 s 11200 75624 12000 75744 6 wbm_a_dat_i[27]
port 57 nsew signal input
rlabel metal3 s 11200 76304 12000 76424 6 wbm_a_dat_i[28]
port 58 nsew signal input
rlabel metal3 s 11200 77120 12000 77240 6 wbm_a_dat_i[29]
port 59 nsew signal input
rlabel metal3 s 11200 56312 12000 56432 6 wbm_a_dat_i[2]
port 60 nsew signal input
rlabel metal3 s 11200 77936 12000 78056 6 wbm_a_dat_i[30]
port 61 nsew signal input
rlabel metal3 s 11200 78616 12000 78736 6 wbm_a_dat_i[31]
port 62 nsew signal input
rlabel metal3 s 11200 57128 12000 57248 6 wbm_a_dat_i[3]
port 63 nsew signal input
rlabel metal3 s 11200 57944 12000 58064 6 wbm_a_dat_i[4]
port 64 nsew signal input
rlabel metal3 s 11200 58624 12000 58744 6 wbm_a_dat_i[5]
port 65 nsew signal input
rlabel metal3 s 11200 59440 12000 59560 6 wbm_a_dat_i[6]
port 66 nsew signal input
rlabel metal3 s 11200 60256 12000 60376 6 wbm_a_dat_i[7]
port 67 nsew signal input
rlabel metal3 s 11200 60936 12000 61056 6 wbm_a_dat_i[8]
port 68 nsew signal input
rlabel metal3 s 11200 61752 12000 61872 6 wbm_a_dat_i[9]
port 69 nsew signal input
rlabel metal3 s 11200 30200 12000 30320 6 wbm_a_dat_o[0]
port 70 nsew signal tristate
rlabel metal3 s 11200 37952 12000 38072 6 wbm_a_dat_o[10]
port 71 nsew signal tristate
rlabel metal3 s 11200 38632 12000 38752 6 wbm_a_dat_o[11]
port 72 nsew signal tristate
rlabel metal3 s 11200 39448 12000 39568 6 wbm_a_dat_o[12]
port 73 nsew signal tristate
rlabel metal3 s 11200 40264 12000 40384 6 wbm_a_dat_o[13]
port 74 nsew signal tristate
rlabel metal3 s 11200 40944 12000 41064 6 wbm_a_dat_o[14]
port 75 nsew signal tristate
rlabel metal3 s 11200 41760 12000 41880 6 wbm_a_dat_o[15]
port 76 nsew signal tristate
rlabel metal3 s 11200 42440 12000 42560 6 wbm_a_dat_o[16]
port 77 nsew signal tristate
rlabel metal3 s 11200 43256 12000 43376 6 wbm_a_dat_o[17]
port 78 nsew signal tristate
rlabel metal3 s 11200 44072 12000 44192 6 wbm_a_dat_o[18]
port 79 nsew signal tristate
rlabel metal3 s 11200 44752 12000 44872 6 wbm_a_dat_o[19]
port 80 nsew signal tristate
rlabel metal3 s 11200 31016 12000 31136 6 wbm_a_dat_o[1]
port 81 nsew signal tristate
rlabel metal3 s 11200 45568 12000 45688 6 wbm_a_dat_o[20]
port 82 nsew signal tristate
rlabel metal3 s 11200 46384 12000 46504 6 wbm_a_dat_o[21]
port 83 nsew signal tristate
rlabel metal3 s 11200 47064 12000 47184 6 wbm_a_dat_o[22]
port 84 nsew signal tristate
rlabel metal3 s 11200 47880 12000 48000 6 wbm_a_dat_o[23]
port 85 nsew signal tristate
rlabel metal3 s 11200 48696 12000 48816 6 wbm_a_dat_o[24]
port 86 nsew signal tristate
rlabel metal3 s 11200 49376 12000 49496 6 wbm_a_dat_o[25]
port 87 nsew signal tristate
rlabel metal3 s 11200 50192 12000 50312 6 wbm_a_dat_o[26]
port 88 nsew signal tristate
rlabel metal3 s 11200 51008 12000 51128 6 wbm_a_dat_o[27]
port 89 nsew signal tristate
rlabel metal3 s 11200 51688 12000 51808 6 wbm_a_dat_o[28]
port 90 nsew signal tristate
rlabel metal3 s 11200 52504 12000 52624 6 wbm_a_dat_o[29]
port 91 nsew signal tristate
rlabel metal3 s 11200 31696 12000 31816 6 wbm_a_dat_o[2]
port 92 nsew signal tristate
rlabel metal3 s 11200 53320 12000 53440 6 wbm_a_dat_o[30]
port 93 nsew signal tristate
rlabel metal3 s 11200 54000 12000 54120 6 wbm_a_dat_o[31]
port 94 nsew signal tristate
rlabel metal3 s 11200 32512 12000 32632 6 wbm_a_dat_o[3]
port 95 nsew signal tristate
rlabel metal3 s 11200 33328 12000 33448 6 wbm_a_dat_o[4]
port 96 nsew signal tristate
rlabel metal3 s 11200 34008 12000 34128 6 wbm_a_dat_o[5]
port 97 nsew signal tristate
rlabel metal3 s 11200 34824 12000 34944 6 wbm_a_dat_o[6]
port 98 nsew signal tristate
rlabel metal3 s 11200 35640 12000 35760 6 wbm_a_dat_o[7]
port 99 nsew signal tristate
rlabel metal3 s 11200 36320 12000 36440 6 wbm_a_dat_o[8]
port 100 nsew signal tristate
rlabel metal3 s 11200 37136 12000 37256 6 wbm_a_dat_o[9]
port 101 nsew signal tristate
rlabel metal3 s 11200 2456 12000 2576 6 wbm_a_sel_o[0]
port 102 nsew signal tristate
rlabel metal3 s 11200 3272 12000 3392 6 wbm_a_sel_o[1]
port 103 nsew signal tristate
rlabel metal3 s 11200 4088 12000 4208 6 wbm_a_sel_o[2]
port 104 nsew signal tristate
rlabel metal3 s 11200 4768 12000 4888 6 wbm_a_sel_o[3]
port 105 nsew signal tristate
rlabel metal3 s 11200 280 12000 400 6 wbm_a_stb_o
port 106 nsew signal tristate
rlabel metal3 s 11200 1776 12000 1896 6 wbm_a_we_o
port 107 nsew signal tristate
rlabel metal3 s 0 79568 800 79688 6 wbm_b_ack_i
port 108 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 wbm_b_adr_o[0]
port 109 nsew signal tristate
rlabel metal3 s 0 48288 800 48408 6 wbm_b_adr_o[1]
port 110 nsew signal tristate
rlabel metal3 s 0 48696 800 48816 6 wbm_b_adr_o[2]
port 111 nsew signal tristate
rlabel metal3 s 0 49104 800 49224 6 wbm_b_adr_o[3]
port 112 nsew signal tristate
rlabel metal3 s 0 49512 800 49632 6 wbm_b_adr_o[4]
port 113 nsew signal tristate
rlabel metal3 s 0 49920 800 50040 6 wbm_b_adr_o[5]
port 114 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 wbm_b_adr_o[6]
port 115 nsew signal tristate
rlabel metal3 s 0 50872 800 50992 6 wbm_b_adr_o[7]
port 116 nsew signal tristate
rlabel metal3 s 0 51280 800 51400 6 wbm_b_adr_o[8]
port 117 nsew signal tristate
rlabel metal3 s 0 51688 800 51808 6 wbm_b_adr_o[9]
port 118 nsew signal tristate
rlabel metal3 s 0 45160 800 45280 6 wbm_b_cyc_o
port 119 nsew signal tristate
rlabel metal3 s 0 65832 800 65952 6 wbm_b_dat_i[0]
port 120 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbm_b_dat_i[10]
port 121 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 wbm_b_dat_i[11]
port 122 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wbm_b_dat_i[12]
port 123 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 wbm_b_dat_i[13]
port 124 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 wbm_b_dat_i[14]
port 125 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbm_b_dat_i[15]
port 126 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wbm_b_dat_i[16]
port 127 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 wbm_b_dat_i[17]
port 128 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 wbm_b_dat_i[18]
port 129 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 wbm_b_dat_i[19]
port 130 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 wbm_b_dat_i[1]
port 131 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 wbm_b_dat_i[20]
port 132 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 wbm_b_dat_i[21]
port 133 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 wbm_b_dat_i[22]
port 134 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 wbm_b_dat_i[23]
port 135 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbm_b_dat_i[24]
port 136 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 wbm_b_dat_i[25]
port 137 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 wbm_b_dat_i[26]
port 138 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wbm_b_dat_i[27]
port 139 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wbm_b_dat_i[28]
port 140 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 wbm_b_dat_i[29]
port 141 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 wbm_b_dat_i[2]
port 142 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 wbm_b_dat_i[30]
port 143 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 wbm_b_dat_i[31]
port 144 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 wbm_b_dat_i[3]
port 145 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 wbm_b_dat_i[4]
port 146 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 wbm_b_dat_i[5]
port 147 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 wbm_b_dat_i[6]
port 148 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 wbm_b_dat_i[7]
port 149 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wbm_b_dat_i[8]
port 150 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 wbm_b_dat_i[9]
port 151 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 wbm_b_dat_o[0]
port 152 nsew signal tristate
rlabel metal3 s 0 56448 800 56568 6 wbm_b_dat_o[10]
port 153 nsew signal tristate
rlabel metal3 s 0 56856 800 56976 6 wbm_b_dat_o[11]
port 154 nsew signal tristate
rlabel metal3 s 0 57264 800 57384 6 wbm_b_dat_o[12]
port 155 nsew signal tristate
rlabel metal3 s 0 57672 800 57792 6 wbm_b_dat_o[13]
port 156 nsew signal tristate
rlabel metal3 s 0 58080 800 58200 6 wbm_b_dat_o[14]
port 157 nsew signal tristate
rlabel metal3 s 0 58488 800 58608 6 wbm_b_dat_o[15]
port 158 nsew signal tristate
rlabel metal3 s 0 59032 800 59152 6 wbm_b_dat_o[16]
port 159 nsew signal tristate
rlabel metal3 s 0 59440 800 59560 6 wbm_b_dat_o[17]
port 160 nsew signal tristate
rlabel metal3 s 0 59848 800 59968 6 wbm_b_dat_o[18]
port 161 nsew signal tristate
rlabel metal3 s 0 60256 800 60376 6 wbm_b_dat_o[19]
port 162 nsew signal tristate
rlabel metal3 s 0 52504 800 52624 6 wbm_b_dat_o[1]
port 163 nsew signal tristate
rlabel metal3 s 0 60664 800 60784 6 wbm_b_dat_o[20]
port 164 nsew signal tristate
rlabel metal3 s 0 61072 800 61192 6 wbm_b_dat_o[21]
port 165 nsew signal tristate
rlabel metal3 s 0 61616 800 61736 6 wbm_b_dat_o[22]
port 166 nsew signal tristate
rlabel metal3 s 0 62024 800 62144 6 wbm_b_dat_o[23]
port 167 nsew signal tristate
rlabel metal3 s 0 62432 800 62552 6 wbm_b_dat_o[24]
port 168 nsew signal tristate
rlabel metal3 s 0 62840 800 62960 6 wbm_b_dat_o[25]
port 169 nsew signal tristate
rlabel metal3 s 0 63248 800 63368 6 wbm_b_dat_o[26]
port 170 nsew signal tristate
rlabel metal3 s 0 63656 800 63776 6 wbm_b_dat_o[27]
port 171 nsew signal tristate
rlabel metal3 s 0 64200 800 64320 6 wbm_b_dat_o[28]
port 172 nsew signal tristate
rlabel metal3 s 0 64608 800 64728 6 wbm_b_dat_o[29]
port 173 nsew signal tristate
rlabel metal3 s 0 52912 800 53032 6 wbm_b_dat_o[2]
port 174 nsew signal tristate
rlabel metal3 s 0 65016 800 65136 6 wbm_b_dat_o[30]
port 175 nsew signal tristate
rlabel metal3 s 0 65424 800 65544 6 wbm_b_dat_o[31]
port 176 nsew signal tristate
rlabel metal3 s 0 53456 800 53576 6 wbm_b_dat_o[3]
port 177 nsew signal tristate
rlabel metal3 s 0 53864 800 53984 6 wbm_b_dat_o[4]
port 178 nsew signal tristate
rlabel metal3 s 0 54272 800 54392 6 wbm_b_dat_o[5]
port 179 nsew signal tristate
rlabel metal3 s 0 54680 800 54800 6 wbm_b_dat_o[6]
port 180 nsew signal tristate
rlabel metal3 s 0 55088 800 55208 6 wbm_b_dat_o[7]
port 181 nsew signal tristate
rlabel metal3 s 0 55496 800 55616 6 wbm_b_dat_o[8]
port 182 nsew signal tristate
rlabel metal3 s 0 55904 800 56024 6 wbm_b_dat_o[9]
port 183 nsew signal tristate
rlabel metal3 s 0 46112 800 46232 6 wbm_b_sel_o[0]
port 184 nsew signal tristate
rlabel metal3 s 0 46520 800 46640 6 wbm_b_sel_o[1]
port 185 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 wbm_b_sel_o[2]
port 186 nsew signal tristate
rlabel metal3 s 0 47336 800 47456 6 wbm_b_sel_o[3]
port 187 nsew signal tristate
rlabel metal3 s 0 44752 800 44872 6 wbm_b_stb_o
port 188 nsew signal tristate
rlabel metal3 s 0 45704 800 45824 6 wbm_b_we_o
port 189 nsew signal tristate
rlabel metal3 s 0 44344 800 44464 6 wbs_ack_o
port 190 nsew signal tristate
rlabel metal3 s 0 3136 800 3256 6 wbs_adr_i[0]
port 191 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wbs_adr_i[10]
port 192 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wbs_adr_i[11]
port 193 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 wbs_adr_i[12]
port 194 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 wbs_adr_i[13]
port 195 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_adr_i[14]
port 196 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_adr_i[15]
port 197 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 wbs_adr_i[16]
port 198 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_adr_i[17]
port 199 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_adr_i[18]
port 200 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 wbs_adr_i[19]
port 201 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 wbs_adr_i[1]
port 202 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 wbs_adr_i[20]
port 203 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 wbs_adr_i[21]
port 204 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 wbs_adr_i[22]
port 205 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_adr_i[23]
port 206 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 wbs_adr_i[24]
port 207 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wbs_adr_i[25]
port 208 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 wbs_adr_i[26]
port 209 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 wbs_adr_i[27]
port 210 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 wbs_adr_i[28]
port 211 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 wbs_adr_i[29]
port 212 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_adr_i[2]
port 213 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 wbs_adr_i[30]
port 214 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wbs_adr_i[31]
port 215 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wbs_adr_i[3]
port 216 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_adr_i[4]
port 217 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wbs_adr_i[5]
port 218 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 wbs_adr_i[6]
port 219 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_adr_i[7]
port 220 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 wbs_adr_i[8]
port 221 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 wbs_adr_i[9]
port 222 nsew signal input
rlabel metal3 s 0 552 800 672 6 wbs_cyc_i
port 223 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wbs_dat_i[0]
port 224 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_i[10]
port 225 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wbs_dat_i[11]
port 226 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 wbs_dat_i[12]
port 227 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wbs_dat_i[13]
port 228 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 wbs_dat_i[14]
port 229 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 wbs_dat_i[15]
port 230 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 wbs_dat_i[16]
port 231 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 wbs_dat_i[17]
port 232 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 wbs_dat_i[18]
port 233 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 wbs_dat_i[19]
port 234 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 wbs_dat_i[1]
port 235 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 wbs_dat_i[20]
port 236 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_i[21]
port 237 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 wbs_dat_i[22]
port 238 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wbs_dat_i[23]
port 239 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wbs_dat_i[24]
port 240 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 wbs_dat_i[25]
port 241 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 wbs_dat_i[26]
port 242 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 wbs_dat_i[27]
port 243 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 wbs_dat_i[28]
port 244 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_i[29]
port 245 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wbs_dat_i[2]
port 246 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 wbs_dat_i[30]
port 247 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 wbs_dat_i[31]
port 248 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wbs_dat_i[3]
port 249 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wbs_dat_i[4]
port 250 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_i[5]
port 251 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wbs_dat_i[6]
port 252 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 wbs_dat_i[7]
port 253 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wbs_dat_i[8]
port 254 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wbs_dat_i[9]
port 255 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 wbs_dat_o[0]
port 256 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_o[10]
port 257 nsew signal tristate
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_o[11]
port 258 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wbs_dat_o[12]
port 259 nsew signal tristate
rlabel metal3 s 0 36184 800 36304 6 wbs_dat_o[13]
port 260 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wbs_dat_o[14]
port 261 nsew signal tristate
rlabel metal3 s 0 37000 800 37120 6 wbs_dat_o[15]
port 262 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wbs_dat_o[16]
port 263 nsew signal tristate
rlabel metal3 s 0 37952 800 38072 6 wbs_dat_o[17]
port 264 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wbs_dat_o[18]
port 265 nsew signal tristate
rlabel metal3 s 0 38768 800 38888 6 wbs_dat_o[19]
port 266 nsew signal tristate
rlabel metal3 s 0 31016 800 31136 6 wbs_dat_o[1]
port 267 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wbs_dat_o[20]
port 268 nsew signal tristate
rlabel metal3 s 0 39584 800 39704 6 wbs_dat_o[21]
port 269 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_o[22]
port 270 nsew signal tristate
rlabel metal3 s 0 40536 800 40656 6 wbs_dat_o[23]
port 271 nsew signal tristate
rlabel metal3 s 0 40944 800 41064 6 wbs_dat_o[24]
port 272 nsew signal tristate
rlabel metal3 s 0 41352 800 41472 6 wbs_dat_o[25]
port 273 nsew signal tristate
rlabel metal3 s 0 41760 800 41880 6 wbs_dat_o[26]
port 274 nsew signal tristate
rlabel metal3 s 0 42168 800 42288 6 wbs_dat_o[27]
port 275 nsew signal tristate
rlabel metal3 s 0 42576 800 42696 6 wbs_dat_o[28]
port 276 nsew signal tristate
rlabel metal3 s 0 43120 800 43240 6 wbs_dat_o[29]
port 277 nsew signal tristate
rlabel metal3 s 0 31424 800 31544 6 wbs_dat_o[2]
port 278 nsew signal tristate
rlabel metal3 s 0 43528 800 43648 6 wbs_dat_o[30]
port 279 nsew signal tristate
rlabel metal3 s 0 43936 800 44056 6 wbs_dat_o[31]
port 280 nsew signal tristate
rlabel metal3 s 0 31832 800 31952 6 wbs_dat_o[3]
port 281 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wbs_dat_o[4]
port 282 nsew signal tristate
rlabel metal3 s 0 32784 800 32904 6 wbs_dat_o[5]
port 283 nsew signal tristate
rlabel metal3 s 0 33192 800 33312 6 wbs_dat_o[6]
port 284 nsew signal tristate
rlabel metal3 s 0 33600 800 33720 6 wbs_dat_o[7]
port 285 nsew signal tristate
rlabel metal3 s 0 34008 800 34128 6 wbs_dat_o[8]
port 286 nsew signal tristate
rlabel metal3 s 0 34416 800 34536 6 wbs_dat_o[9]
port 287 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wbs_sel_i[0]
port 288 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 wbs_sel_i[1]
port 289 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wbs_sel_i[2]
port 290 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wbs_sel_i[3]
port 291 nsew signal input
rlabel metal3 s 0 144 800 264 6 wbs_stb_i
port 292 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_we_i
port 293 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
