VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_bridge_2way
  CLASS BLOCK ;
  FOREIGN wb_bridge_2way ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 400.000 ;
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 12.875 10.640 14.475 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.195 10.640 30.795 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.515 10.640 47.115 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.035 10.640 22.635 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.355 10.640 38.955 389.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 397.160 60.000 397.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END wb_rst_i
  PIN wbm_a_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 393.080 60.000 393.680 ;
    END
  END wbm_a_ack_i
  PIN wbm_a_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 27.920 60.000 28.520 ;
    END
  END wbm_a_adr_o[0]
  PIN wbm_a_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 66.000 60.000 66.600 ;
    END
  END wbm_a_adr_o[10]
  PIN wbm_a_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 69.400 60.000 70.000 ;
    END
  END wbm_a_adr_o[11]
  PIN wbm_a_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 73.480 60.000 74.080 ;
    END
  END wbm_a_adr_o[12]
  PIN wbm_a_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 77.560 60.000 78.160 ;
    END
  END wbm_a_adr_o[13]
  PIN wbm_a_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 80.960 60.000 81.560 ;
    END
  END wbm_a_adr_o[14]
  PIN wbm_a_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 85.040 60.000 85.640 ;
    END
  END wbm_a_adr_o[15]
  PIN wbm_a_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 88.440 60.000 89.040 ;
    END
  END wbm_a_adr_o[16]
  PIN wbm_a_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 92.520 60.000 93.120 ;
    END
  END wbm_a_adr_o[17]
  PIN wbm_a_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 96.600 60.000 97.200 ;
    END
  END wbm_a_adr_o[18]
  PIN wbm_a_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 100.000 60.000 100.600 ;
    END
  END wbm_a_adr_o[19]
  PIN wbm_a_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 31.320 60.000 31.920 ;
    END
  END wbm_a_adr_o[1]
  PIN wbm_a_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 104.080 60.000 104.680 ;
    END
  END wbm_a_adr_o[20]
  PIN wbm_a_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 107.480 60.000 108.080 ;
    END
  END wbm_a_adr_o[21]
  PIN wbm_a_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 111.560 60.000 112.160 ;
    END
  END wbm_a_adr_o[22]
  PIN wbm_a_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 115.640 60.000 116.240 ;
    END
  END wbm_a_adr_o[23]
  PIN wbm_a_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 119.040 60.000 119.640 ;
    END
  END wbm_a_adr_o[24]
  PIN wbm_a_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 123.120 60.000 123.720 ;
    END
  END wbm_a_adr_o[25]
  PIN wbm_a_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 126.520 60.000 127.120 ;
    END
  END wbm_a_adr_o[26]
  PIN wbm_a_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 130.600 60.000 131.200 ;
    END
  END wbm_a_adr_o[27]
  PIN wbm_a_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 134.680 60.000 135.280 ;
    END
  END wbm_a_adr_o[28]
  PIN wbm_a_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 138.080 60.000 138.680 ;
    END
  END wbm_a_adr_o[29]
  PIN wbm_a_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 35.400 60.000 36.000 ;
    END
  END wbm_a_adr_o[2]
  PIN wbm_a_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 142.160 60.000 142.760 ;
    END
  END wbm_a_adr_o[30]
  PIN wbm_a_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 145.560 60.000 146.160 ;
    END
  END wbm_a_adr_o[31]
  PIN wbm_a_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 39.480 60.000 40.080 ;
    END
  END wbm_a_adr_o[3]
  PIN wbm_a_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 42.880 60.000 43.480 ;
    END
  END wbm_a_adr_o[4]
  PIN wbm_a_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 46.960 60.000 47.560 ;
    END
  END wbm_a_adr_o[5]
  PIN wbm_a_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 50.360 60.000 50.960 ;
    END
  END wbm_a_adr_o[6]
  PIN wbm_a_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 54.440 60.000 55.040 ;
    END
  END wbm_a_adr_o[7]
  PIN wbm_a_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 58.520 60.000 59.120 ;
    END
  END wbm_a_adr_o[8]
  PIN wbm_a_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 61.920 60.000 62.520 ;
    END
  END wbm_a_adr_o[9]
  PIN wbm_a_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 4.800 60.000 5.400 ;
    END
  END wbm_a_cyc_o
  PIN wbm_a_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 271.360 60.000 271.960 ;
    END
  END wbm_a_dat_i[0]
  PIN wbm_a_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 309.440 60.000 310.040 ;
    END
  END wbm_a_dat_i[10]
  PIN wbm_a_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 313.520 60.000 314.120 ;
    END
  END wbm_a_dat_i[11]
  PIN wbm_a_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 316.920 60.000 317.520 ;
    END
  END wbm_a_dat_i[12]
  PIN wbm_a_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 321.000 60.000 321.600 ;
    END
  END wbm_a_dat_i[13]
  PIN wbm_a_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 325.080 60.000 325.680 ;
    END
  END wbm_a_dat_i[14]
  PIN wbm_a_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 328.480 60.000 329.080 ;
    END
  END wbm_a_dat_i[15]
  PIN wbm_a_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 332.560 60.000 333.160 ;
    END
  END wbm_a_dat_i[16]
  PIN wbm_a_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 335.960 60.000 336.560 ;
    END
  END wbm_a_dat_i[17]
  PIN wbm_a_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 340.040 60.000 340.640 ;
    END
  END wbm_a_dat_i[18]
  PIN wbm_a_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 344.120 60.000 344.720 ;
    END
  END wbm_a_dat_i[19]
  PIN wbm_a_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 275.440 60.000 276.040 ;
    END
  END wbm_a_dat_i[1]
  PIN wbm_a_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 347.520 60.000 348.120 ;
    END
  END wbm_a_dat_i[20]
  PIN wbm_a_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 351.600 60.000 352.200 ;
    END
  END wbm_a_dat_i[21]
  PIN wbm_a_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 355.000 60.000 355.600 ;
    END
  END wbm_a_dat_i[22]
  PIN wbm_a_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 359.080 60.000 359.680 ;
    END
  END wbm_a_dat_i[23]
  PIN wbm_a_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 363.160 60.000 363.760 ;
    END
  END wbm_a_dat_i[24]
  PIN wbm_a_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 366.560 60.000 367.160 ;
    END
  END wbm_a_dat_i[25]
  PIN wbm_a_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 370.640 60.000 371.240 ;
    END
  END wbm_a_dat_i[26]
  PIN wbm_a_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 374.040 60.000 374.640 ;
    END
  END wbm_a_dat_i[27]
  PIN wbm_a_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 378.120 60.000 378.720 ;
    END
  END wbm_a_dat_i[28]
  PIN wbm_a_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 382.200 60.000 382.800 ;
    END
  END wbm_a_dat_i[29]
  PIN wbm_a_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 278.840 60.000 279.440 ;
    END
  END wbm_a_dat_i[2]
  PIN wbm_a_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 385.600 60.000 386.200 ;
    END
  END wbm_a_dat_i[30]
  PIN wbm_a_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 389.680 60.000 390.280 ;
    END
  END wbm_a_dat_i[31]
  PIN wbm_a_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 282.920 60.000 283.520 ;
    END
  END wbm_a_dat_i[3]
  PIN wbm_a_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 287.000 60.000 287.600 ;
    END
  END wbm_a_dat_i[4]
  PIN wbm_a_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 290.400 60.000 291.000 ;
    END
  END wbm_a_dat_i[5]
  PIN wbm_a_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 294.480 60.000 295.080 ;
    END
  END wbm_a_dat_i[6]
  PIN wbm_a_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 297.880 60.000 298.480 ;
    END
  END wbm_a_dat_i[7]
  PIN wbm_a_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 301.960 60.000 302.560 ;
    END
  END wbm_a_dat_i[8]
  PIN wbm_a_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 306.040 60.000 306.640 ;
    END
  END wbm_a_dat_i[9]
  PIN wbm_a_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 149.640 60.000 150.240 ;
    END
  END wbm_a_dat_o[0]
  PIN wbm_a_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 187.720 60.000 188.320 ;
    END
  END wbm_a_dat_o[10]
  PIN wbm_a_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 191.800 60.000 192.400 ;
    END
  END wbm_a_dat_o[11]
  PIN wbm_a_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 195.200 60.000 195.800 ;
    END
  END wbm_a_dat_o[12]
  PIN wbm_a_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 199.280 60.000 199.880 ;
    END
  END wbm_a_dat_o[13]
  PIN wbm_a_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 202.680 60.000 203.280 ;
    END
  END wbm_a_dat_o[14]
  PIN wbm_a_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 206.760 60.000 207.360 ;
    END
  END wbm_a_dat_o[15]
  PIN wbm_a_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 210.840 60.000 211.440 ;
    END
  END wbm_a_dat_o[16]
  PIN wbm_a_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 214.240 60.000 214.840 ;
    END
  END wbm_a_dat_o[17]
  PIN wbm_a_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 218.320 60.000 218.920 ;
    END
  END wbm_a_dat_o[18]
  PIN wbm_a_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 221.720 60.000 222.320 ;
    END
  END wbm_a_dat_o[19]
  PIN wbm_a_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 153.720 60.000 154.320 ;
    END
  END wbm_a_dat_o[1]
  PIN wbm_a_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 225.800 60.000 226.400 ;
    END
  END wbm_a_dat_o[20]
  PIN wbm_a_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 229.880 60.000 230.480 ;
    END
  END wbm_a_dat_o[21]
  PIN wbm_a_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 233.280 60.000 233.880 ;
    END
  END wbm_a_dat_o[22]
  PIN wbm_a_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 237.360 60.000 237.960 ;
    END
  END wbm_a_dat_o[23]
  PIN wbm_a_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 240.760 60.000 241.360 ;
    END
  END wbm_a_dat_o[24]
  PIN wbm_a_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 244.840 60.000 245.440 ;
    END
  END wbm_a_dat_o[25]
  PIN wbm_a_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 248.920 60.000 249.520 ;
    END
  END wbm_a_dat_o[26]
  PIN wbm_a_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 252.320 60.000 252.920 ;
    END
  END wbm_a_dat_o[27]
  PIN wbm_a_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 256.400 60.000 257.000 ;
    END
  END wbm_a_dat_o[28]
  PIN wbm_a_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 259.800 60.000 260.400 ;
    END
  END wbm_a_dat_o[29]
  PIN wbm_a_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 157.120 60.000 157.720 ;
    END
  END wbm_a_dat_o[2]
  PIN wbm_a_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 263.880 60.000 264.480 ;
    END
  END wbm_a_dat_o[30]
  PIN wbm_a_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 267.960 60.000 268.560 ;
    END
  END wbm_a_dat_o[31]
  PIN wbm_a_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 161.200 60.000 161.800 ;
    END
  END wbm_a_dat_o[3]
  PIN wbm_a_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 164.600 60.000 165.200 ;
    END
  END wbm_a_dat_o[4]
  PIN wbm_a_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 168.680 60.000 169.280 ;
    END
  END wbm_a_dat_o[5]
  PIN wbm_a_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 172.760 60.000 173.360 ;
    END
  END wbm_a_dat_o[6]
  PIN wbm_a_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 176.160 60.000 176.760 ;
    END
  END wbm_a_dat_o[7]
  PIN wbm_a_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 180.240 60.000 180.840 ;
    END
  END wbm_a_dat_o[8]
  PIN wbm_a_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 183.640 60.000 184.240 ;
    END
  END wbm_a_dat_o[9]
  PIN wbm_a_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 12.280 60.000 12.880 ;
    END
  END wbm_a_sel_o[0]
  PIN wbm_a_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 16.360 60.000 16.960 ;
    END
  END wbm_a_sel_o[1]
  PIN wbm_a_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 20.440 60.000 21.040 ;
    END
  END wbm_a_sel_o[2]
  PIN wbm_a_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 23.840 60.000 24.440 ;
    END
  END wbm_a_sel_o[3]
  PIN wbm_a_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 1.400 60.000 2.000 ;
    END
  END wbm_a_stb_o
  PIN wbm_a_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 56.000 8.880 60.000 9.480 ;
    END
  END wbm_a_we_o
  PIN wbm_b_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END wbm_b_ack_i
  PIN wbm_b_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END wbm_b_adr_o[0]
  PIN wbm_b_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END wbm_b_adr_o[1]
  PIN wbm_b_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END wbm_b_adr_o[2]
  PIN wbm_b_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END wbm_b_adr_o[3]
  PIN wbm_b_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END wbm_b_adr_o[4]
  PIN wbm_b_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END wbm_b_adr_o[5]
  PIN wbm_b_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END wbm_b_adr_o[6]
  PIN wbm_b_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END wbm_b_adr_o[7]
  PIN wbm_b_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END wbm_b_adr_o[8]
  PIN wbm_b_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END wbm_b_adr_o[9]
  PIN wbm_b_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END wbm_b_cyc_o
  PIN wbm_b_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wbm_b_dat_i[0]
  PIN wbm_b_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wbm_b_dat_i[10]
  PIN wbm_b_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END wbm_b_dat_i[11]
  PIN wbm_b_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END wbm_b_dat_i[12]
  PIN wbm_b_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END wbm_b_dat_i[13]
  PIN wbm_b_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END wbm_b_dat_i[14]
  PIN wbm_b_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wbm_b_dat_i[15]
  PIN wbm_b_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END wbm_b_dat_i[16]
  PIN wbm_b_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END wbm_b_dat_i[17]
  PIN wbm_b_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.920 4.000 368.520 ;
    END
  END wbm_b_dat_i[18]
  PIN wbm_b_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END wbm_b_dat_i[19]
  PIN wbm_b_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END wbm_b_dat_i[1]
  PIN wbm_b_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END wbm_b_dat_i[20]
  PIN wbm_b_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END wbm_b_dat_i[21]
  PIN wbm_b_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END wbm_b_dat_i[22]
  PIN wbm_b_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END wbm_b_dat_i[23]
  PIN wbm_b_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wbm_b_dat_i[24]
  PIN wbm_b_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END wbm_b_dat_i[25]
  PIN wbm_b_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END wbm_b_dat_i[26]
  PIN wbm_b_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wbm_b_dat_i[27]
  PIN wbm_b_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END wbm_b_dat_i[28]
  PIN wbm_b_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END wbm_b_dat_i[29]
  PIN wbm_b_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END wbm_b_dat_i[2]
  PIN wbm_b_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END wbm_b_dat_i[30]
  PIN wbm_b_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END wbm_b_dat_i[31]
  PIN wbm_b_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END wbm_b_dat_i[3]
  PIN wbm_b_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END wbm_b_dat_i[4]
  PIN wbm_b_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END wbm_b_dat_i[5]
  PIN wbm_b_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END wbm_b_dat_i[6]
  PIN wbm_b_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END wbm_b_dat_i[7]
  PIN wbm_b_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END wbm_b_dat_i[8]
  PIN wbm_b_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END wbm_b_dat_i[9]
  PIN wbm_b_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END wbm_b_dat_o[0]
  PIN wbm_b_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END wbm_b_dat_o[10]
  PIN wbm_b_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END wbm_b_dat_o[11]
  PIN wbm_b_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END wbm_b_dat_o[12]
  PIN wbm_b_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END wbm_b_dat_o[13]
  PIN wbm_b_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END wbm_b_dat_o[14]
  PIN wbm_b_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END wbm_b_dat_o[15]
  PIN wbm_b_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END wbm_b_dat_o[16]
  PIN wbm_b_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END wbm_b_dat_o[17]
  PIN wbm_b_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END wbm_b_dat_o[18]
  PIN wbm_b_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.280 4.000 301.880 ;
    END
  END wbm_b_dat_o[19]
  PIN wbm_b_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END wbm_b_dat_o[1]
  PIN wbm_b_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END wbm_b_dat_o[20]
  PIN wbm_b_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 305.360 4.000 305.960 ;
    END
  END wbm_b_dat_o[21]
  PIN wbm_b_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END wbm_b_dat_o[22]
  PIN wbm_b_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END wbm_b_dat_o[23]
  PIN wbm_b_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END wbm_b_dat_o[24]
  PIN wbm_b_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END wbm_b_dat_o[25]
  PIN wbm_b_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END wbm_b_dat_o[26]
  PIN wbm_b_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wbm_b_dat_o[27]
  PIN wbm_b_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END wbm_b_dat_o[28]
  PIN wbm_b_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wbm_b_dat_o[29]
  PIN wbm_b_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END wbm_b_dat_o[2]
  PIN wbm_b_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END wbm_b_dat_o[30]
  PIN wbm_b_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END wbm_b_dat_o[31]
  PIN wbm_b_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END wbm_b_dat_o[3]
  PIN wbm_b_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END wbm_b_dat_o[4]
  PIN wbm_b_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END wbm_b_dat_o[5]
  PIN wbm_b_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END wbm_b_dat_o[6]
  PIN wbm_b_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END wbm_b_dat_o[7]
  PIN wbm_b_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END wbm_b_dat_o[8]
  PIN wbm_b_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END wbm_b_dat_o[9]
  PIN wbm_b_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END wbm_b_sel_o[0]
  PIN wbm_b_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END wbm_b_sel_o[1]
  PIN wbm_b_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END wbm_b_sel_o[2]
  PIN wbm_b_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END wbm_b_sel_o[3]
  PIN wbm_b_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END wbm_b_stb_o
  PIN wbm_b_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END wbm_b_we_o
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.960 4.000 183.560 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.920 4.000 198.520 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.080 4.000 172.680 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 3.825 10.795 59.655 389.895 ;
      LAYER met1 ;
        RECT 0.530 2.420 59.715 389.940 ;
      LAYER met2 ;
        RECT 0.560 4.280 55.110 398.325 ;
        RECT 0.560 0.835 29.710 4.280 ;
        RECT 30.550 0.835 55.110 4.280 ;
      LAYER met3 ;
        RECT 4.400 398.160 56.000 398.305 ;
        RECT 4.400 397.440 55.600 398.160 ;
        RECT 3.990 396.800 55.600 397.440 ;
        RECT 4.400 396.760 55.600 396.800 ;
        RECT 4.400 395.400 56.000 396.760 ;
        RECT 3.990 394.760 56.000 395.400 ;
        RECT 4.400 394.080 56.000 394.760 ;
        RECT 4.400 393.360 55.600 394.080 ;
        RECT 3.990 392.720 55.600 393.360 ;
        RECT 4.400 392.680 55.600 392.720 ;
        RECT 4.400 391.320 56.000 392.680 ;
        RECT 3.990 390.680 56.000 391.320 ;
        RECT 4.400 389.280 55.600 390.680 ;
        RECT 3.990 388.640 56.000 389.280 ;
        RECT 4.400 387.240 56.000 388.640 ;
        RECT 3.990 386.600 56.000 387.240 ;
        RECT 3.990 385.920 55.600 386.600 ;
        RECT 4.400 385.200 55.600 385.920 ;
        RECT 4.400 384.520 56.000 385.200 ;
        RECT 3.990 383.880 56.000 384.520 ;
        RECT 4.400 383.200 56.000 383.880 ;
        RECT 4.400 382.480 55.600 383.200 ;
        RECT 3.990 381.840 55.600 382.480 ;
        RECT 4.400 381.800 55.600 381.840 ;
        RECT 4.400 380.440 56.000 381.800 ;
        RECT 3.990 379.800 56.000 380.440 ;
        RECT 4.400 379.120 56.000 379.800 ;
        RECT 4.400 378.400 55.600 379.120 ;
        RECT 3.990 377.760 55.600 378.400 ;
        RECT 4.400 377.720 55.600 377.760 ;
        RECT 4.400 376.360 56.000 377.720 ;
        RECT 3.990 375.720 56.000 376.360 ;
        RECT 4.400 375.040 56.000 375.720 ;
        RECT 4.400 374.320 55.600 375.040 ;
        RECT 3.990 373.640 55.600 374.320 ;
        RECT 3.990 373.000 56.000 373.640 ;
        RECT 4.400 371.640 56.000 373.000 ;
        RECT 4.400 371.600 55.600 371.640 ;
        RECT 3.990 370.960 55.600 371.600 ;
        RECT 4.400 370.240 55.600 370.960 ;
        RECT 4.400 369.560 56.000 370.240 ;
        RECT 3.990 368.920 56.000 369.560 ;
        RECT 4.400 367.560 56.000 368.920 ;
        RECT 4.400 367.520 55.600 367.560 ;
        RECT 3.990 366.880 55.600 367.520 ;
        RECT 4.400 366.160 55.600 366.880 ;
        RECT 4.400 365.480 56.000 366.160 ;
        RECT 3.990 364.840 56.000 365.480 ;
        RECT 4.400 364.160 56.000 364.840 ;
        RECT 4.400 363.440 55.600 364.160 ;
        RECT 3.990 362.800 55.600 363.440 ;
        RECT 4.400 362.760 55.600 362.800 ;
        RECT 4.400 361.400 56.000 362.760 ;
        RECT 3.990 360.080 56.000 361.400 ;
        RECT 4.400 358.680 55.600 360.080 ;
        RECT 3.990 358.040 56.000 358.680 ;
        RECT 4.400 356.640 56.000 358.040 ;
        RECT 3.990 356.000 56.000 356.640 ;
        RECT 4.400 354.600 55.600 356.000 ;
        RECT 3.990 353.960 56.000 354.600 ;
        RECT 4.400 352.600 56.000 353.960 ;
        RECT 4.400 352.560 55.600 352.600 ;
        RECT 3.990 351.920 55.600 352.560 ;
        RECT 4.400 351.200 55.600 351.920 ;
        RECT 4.400 350.520 56.000 351.200 ;
        RECT 3.990 349.880 56.000 350.520 ;
        RECT 4.400 348.520 56.000 349.880 ;
        RECT 4.400 348.480 55.600 348.520 ;
        RECT 3.990 347.160 55.600 348.480 ;
        RECT 4.400 347.120 55.600 347.160 ;
        RECT 4.400 345.760 56.000 347.120 ;
        RECT 3.990 345.120 56.000 345.760 ;
        RECT 4.400 343.720 55.600 345.120 ;
        RECT 3.990 343.080 56.000 343.720 ;
        RECT 4.400 341.680 56.000 343.080 ;
        RECT 3.990 341.040 56.000 341.680 ;
        RECT 4.400 339.640 55.600 341.040 ;
        RECT 3.990 339.000 56.000 339.640 ;
        RECT 4.400 337.600 56.000 339.000 ;
        RECT 3.990 336.960 56.000 337.600 ;
        RECT 4.400 335.560 55.600 336.960 ;
        RECT 3.990 334.920 56.000 335.560 ;
        RECT 4.400 333.560 56.000 334.920 ;
        RECT 4.400 333.520 55.600 333.560 ;
        RECT 3.990 332.200 55.600 333.520 ;
        RECT 4.400 332.160 55.600 332.200 ;
        RECT 4.400 330.800 56.000 332.160 ;
        RECT 3.990 330.160 56.000 330.800 ;
        RECT 4.400 329.480 56.000 330.160 ;
        RECT 4.400 328.760 55.600 329.480 ;
        RECT 3.990 328.120 55.600 328.760 ;
        RECT 4.400 328.080 55.600 328.120 ;
        RECT 4.400 326.720 56.000 328.080 ;
        RECT 3.990 326.080 56.000 326.720 ;
        RECT 4.400 324.680 55.600 326.080 ;
        RECT 3.990 324.040 56.000 324.680 ;
        RECT 4.400 322.640 56.000 324.040 ;
        RECT 3.990 322.000 56.000 322.640 ;
        RECT 4.400 320.600 55.600 322.000 ;
        RECT 3.990 319.280 56.000 320.600 ;
        RECT 4.400 317.920 56.000 319.280 ;
        RECT 4.400 317.880 55.600 317.920 ;
        RECT 3.990 317.240 55.600 317.880 ;
        RECT 4.400 316.520 55.600 317.240 ;
        RECT 4.400 315.840 56.000 316.520 ;
        RECT 3.990 315.200 56.000 315.840 ;
        RECT 4.400 314.520 56.000 315.200 ;
        RECT 4.400 313.800 55.600 314.520 ;
        RECT 3.990 313.160 55.600 313.800 ;
        RECT 4.400 313.120 55.600 313.160 ;
        RECT 4.400 311.760 56.000 313.120 ;
        RECT 3.990 311.120 56.000 311.760 ;
        RECT 4.400 310.440 56.000 311.120 ;
        RECT 4.400 309.720 55.600 310.440 ;
        RECT 3.990 309.080 55.600 309.720 ;
        RECT 4.400 309.040 55.600 309.080 ;
        RECT 4.400 307.680 56.000 309.040 ;
        RECT 3.990 307.040 56.000 307.680 ;
        RECT 3.990 306.360 55.600 307.040 ;
        RECT 4.400 305.640 55.600 306.360 ;
        RECT 4.400 304.960 56.000 305.640 ;
        RECT 3.990 304.320 56.000 304.960 ;
        RECT 4.400 302.960 56.000 304.320 ;
        RECT 4.400 302.920 55.600 302.960 ;
        RECT 3.990 302.280 55.600 302.920 ;
        RECT 4.400 301.560 55.600 302.280 ;
        RECT 4.400 300.880 56.000 301.560 ;
        RECT 3.990 300.240 56.000 300.880 ;
        RECT 4.400 298.880 56.000 300.240 ;
        RECT 4.400 298.840 55.600 298.880 ;
        RECT 3.990 298.200 55.600 298.840 ;
        RECT 4.400 297.480 55.600 298.200 ;
        RECT 4.400 296.800 56.000 297.480 ;
        RECT 3.990 296.160 56.000 296.800 ;
        RECT 4.400 295.480 56.000 296.160 ;
        RECT 4.400 294.760 55.600 295.480 ;
        RECT 3.990 294.080 55.600 294.760 ;
        RECT 3.990 293.440 56.000 294.080 ;
        RECT 4.400 292.040 56.000 293.440 ;
        RECT 3.990 291.400 56.000 292.040 ;
        RECT 4.400 290.000 55.600 291.400 ;
        RECT 3.990 289.360 56.000 290.000 ;
        RECT 4.400 288.000 56.000 289.360 ;
        RECT 4.400 287.960 55.600 288.000 ;
        RECT 3.990 287.320 55.600 287.960 ;
        RECT 4.400 286.600 55.600 287.320 ;
        RECT 4.400 285.920 56.000 286.600 ;
        RECT 3.990 285.280 56.000 285.920 ;
        RECT 4.400 283.920 56.000 285.280 ;
        RECT 4.400 283.880 55.600 283.920 ;
        RECT 3.990 283.240 55.600 283.880 ;
        RECT 4.400 282.520 55.600 283.240 ;
        RECT 4.400 281.840 56.000 282.520 ;
        RECT 3.990 280.520 56.000 281.840 ;
        RECT 4.400 279.840 56.000 280.520 ;
        RECT 4.400 279.120 55.600 279.840 ;
        RECT 3.990 278.480 55.600 279.120 ;
        RECT 4.400 278.440 55.600 278.480 ;
        RECT 4.400 277.080 56.000 278.440 ;
        RECT 3.990 276.440 56.000 277.080 ;
        RECT 4.400 275.040 55.600 276.440 ;
        RECT 3.990 274.400 56.000 275.040 ;
        RECT 4.400 273.000 56.000 274.400 ;
        RECT 3.990 272.360 56.000 273.000 ;
        RECT 4.400 270.960 55.600 272.360 ;
        RECT 3.990 270.320 56.000 270.960 ;
        RECT 4.400 268.960 56.000 270.320 ;
        RECT 4.400 268.920 55.600 268.960 ;
        RECT 3.990 268.280 55.600 268.920 ;
        RECT 4.400 267.560 55.600 268.280 ;
        RECT 4.400 266.880 56.000 267.560 ;
        RECT 3.990 265.560 56.000 266.880 ;
        RECT 4.400 264.880 56.000 265.560 ;
        RECT 4.400 264.160 55.600 264.880 ;
        RECT 3.990 263.520 55.600 264.160 ;
        RECT 4.400 263.480 55.600 263.520 ;
        RECT 4.400 262.120 56.000 263.480 ;
        RECT 3.990 261.480 56.000 262.120 ;
        RECT 4.400 260.800 56.000 261.480 ;
        RECT 4.400 260.080 55.600 260.800 ;
        RECT 3.990 259.440 55.600 260.080 ;
        RECT 4.400 259.400 55.600 259.440 ;
        RECT 4.400 258.040 56.000 259.400 ;
        RECT 3.990 257.400 56.000 258.040 ;
        RECT 4.400 256.000 55.600 257.400 ;
        RECT 3.990 255.360 56.000 256.000 ;
        RECT 4.400 253.960 56.000 255.360 ;
        RECT 3.990 253.320 56.000 253.960 ;
        RECT 3.990 252.640 55.600 253.320 ;
        RECT 4.400 251.920 55.600 252.640 ;
        RECT 4.400 251.240 56.000 251.920 ;
        RECT 3.990 250.600 56.000 251.240 ;
        RECT 4.400 249.920 56.000 250.600 ;
        RECT 4.400 249.200 55.600 249.920 ;
        RECT 3.990 248.560 55.600 249.200 ;
        RECT 4.400 248.520 55.600 248.560 ;
        RECT 4.400 247.160 56.000 248.520 ;
        RECT 3.990 246.520 56.000 247.160 ;
        RECT 4.400 245.840 56.000 246.520 ;
        RECT 4.400 245.120 55.600 245.840 ;
        RECT 3.990 244.480 55.600 245.120 ;
        RECT 4.400 244.440 55.600 244.480 ;
        RECT 4.400 243.080 56.000 244.440 ;
        RECT 3.990 242.440 56.000 243.080 ;
        RECT 4.400 241.760 56.000 242.440 ;
        RECT 4.400 241.040 55.600 241.760 ;
        RECT 3.990 240.360 55.600 241.040 ;
        RECT 3.990 239.720 56.000 240.360 ;
        RECT 4.400 238.360 56.000 239.720 ;
        RECT 4.400 238.320 55.600 238.360 ;
        RECT 3.990 237.680 55.600 238.320 ;
        RECT 4.400 236.960 55.600 237.680 ;
        RECT 4.400 236.280 56.000 236.960 ;
        RECT 3.990 235.640 56.000 236.280 ;
        RECT 4.400 234.280 56.000 235.640 ;
        RECT 4.400 234.240 55.600 234.280 ;
        RECT 3.990 233.600 55.600 234.240 ;
        RECT 4.400 232.880 55.600 233.600 ;
        RECT 4.400 232.200 56.000 232.880 ;
        RECT 3.990 231.560 56.000 232.200 ;
        RECT 4.400 230.880 56.000 231.560 ;
        RECT 4.400 230.160 55.600 230.880 ;
        RECT 3.990 229.520 55.600 230.160 ;
        RECT 4.400 229.480 55.600 229.520 ;
        RECT 4.400 228.120 56.000 229.480 ;
        RECT 3.990 226.800 56.000 228.120 ;
        RECT 4.400 225.400 55.600 226.800 ;
        RECT 3.990 224.760 56.000 225.400 ;
        RECT 4.400 223.360 56.000 224.760 ;
        RECT 3.990 222.720 56.000 223.360 ;
        RECT 4.400 221.320 55.600 222.720 ;
        RECT 3.990 220.680 56.000 221.320 ;
        RECT 4.400 219.320 56.000 220.680 ;
        RECT 4.400 219.280 55.600 219.320 ;
        RECT 3.990 218.640 55.600 219.280 ;
        RECT 4.400 217.920 55.600 218.640 ;
        RECT 4.400 217.240 56.000 217.920 ;
        RECT 3.990 216.600 56.000 217.240 ;
        RECT 4.400 215.240 56.000 216.600 ;
        RECT 4.400 215.200 55.600 215.240 ;
        RECT 3.990 213.880 55.600 215.200 ;
        RECT 4.400 213.840 55.600 213.880 ;
        RECT 4.400 212.480 56.000 213.840 ;
        RECT 3.990 211.840 56.000 212.480 ;
        RECT 4.400 210.440 55.600 211.840 ;
        RECT 3.990 209.800 56.000 210.440 ;
        RECT 4.400 208.400 56.000 209.800 ;
        RECT 3.990 207.760 56.000 208.400 ;
        RECT 4.400 206.360 55.600 207.760 ;
        RECT 3.990 205.720 56.000 206.360 ;
        RECT 4.400 204.320 56.000 205.720 ;
        RECT 3.990 203.680 56.000 204.320 ;
        RECT 4.400 202.280 55.600 203.680 ;
        RECT 3.990 201.640 56.000 202.280 ;
        RECT 4.400 200.280 56.000 201.640 ;
        RECT 4.400 200.240 55.600 200.280 ;
        RECT 3.990 198.920 55.600 200.240 ;
        RECT 4.400 198.880 55.600 198.920 ;
        RECT 4.400 197.520 56.000 198.880 ;
        RECT 3.990 196.880 56.000 197.520 ;
        RECT 4.400 196.200 56.000 196.880 ;
        RECT 4.400 195.480 55.600 196.200 ;
        RECT 3.990 194.840 55.600 195.480 ;
        RECT 4.400 194.800 55.600 194.840 ;
        RECT 4.400 193.440 56.000 194.800 ;
        RECT 3.990 192.800 56.000 193.440 ;
        RECT 4.400 191.400 55.600 192.800 ;
        RECT 3.990 190.760 56.000 191.400 ;
        RECT 4.400 189.360 56.000 190.760 ;
        RECT 3.990 188.720 56.000 189.360 ;
        RECT 4.400 187.320 55.600 188.720 ;
        RECT 3.990 186.000 56.000 187.320 ;
        RECT 4.400 184.640 56.000 186.000 ;
        RECT 4.400 184.600 55.600 184.640 ;
        RECT 3.990 183.960 55.600 184.600 ;
        RECT 4.400 183.240 55.600 183.960 ;
        RECT 4.400 182.560 56.000 183.240 ;
        RECT 3.990 181.920 56.000 182.560 ;
        RECT 4.400 181.240 56.000 181.920 ;
        RECT 4.400 180.520 55.600 181.240 ;
        RECT 3.990 179.880 55.600 180.520 ;
        RECT 4.400 179.840 55.600 179.880 ;
        RECT 4.400 178.480 56.000 179.840 ;
        RECT 3.990 177.840 56.000 178.480 ;
        RECT 4.400 177.160 56.000 177.840 ;
        RECT 4.400 176.440 55.600 177.160 ;
        RECT 3.990 175.800 55.600 176.440 ;
        RECT 4.400 175.760 55.600 175.800 ;
        RECT 4.400 174.400 56.000 175.760 ;
        RECT 3.990 173.760 56.000 174.400 ;
        RECT 3.990 173.080 55.600 173.760 ;
        RECT 4.400 172.360 55.600 173.080 ;
        RECT 4.400 171.680 56.000 172.360 ;
        RECT 3.990 171.040 56.000 171.680 ;
        RECT 4.400 169.680 56.000 171.040 ;
        RECT 4.400 169.640 55.600 169.680 ;
        RECT 3.990 169.000 55.600 169.640 ;
        RECT 4.400 168.280 55.600 169.000 ;
        RECT 4.400 167.600 56.000 168.280 ;
        RECT 3.990 166.960 56.000 167.600 ;
        RECT 4.400 165.600 56.000 166.960 ;
        RECT 4.400 165.560 55.600 165.600 ;
        RECT 3.990 164.920 55.600 165.560 ;
        RECT 4.400 164.200 55.600 164.920 ;
        RECT 4.400 163.520 56.000 164.200 ;
        RECT 3.990 162.880 56.000 163.520 ;
        RECT 4.400 162.200 56.000 162.880 ;
        RECT 4.400 161.480 55.600 162.200 ;
        RECT 3.990 160.800 55.600 161.480 ;
        RECT 3.990 160.160 56.000 160.800 ;
        RECT 4.400 158.760 56.000 160.160 ;
        RECT 3.990 158.120 56.000 158.760 ;
        RECT 4.400 156.720 55.600 158.120 ;
        RECT 3.990 156.080 56.000 156.720 ;
        RECT 4.400 154.720 56.000 156.080 ;
        RECT 4.400 154.680 55.600 154.720 ;
        RECT 3.990 154.040 55.600 154.680 ;
        RECT 4.400 153.320 55.600 154.040 ;
        RECT 4.400 152.640 56.000 153.320 ;
        RECT 3.990 152.000 56.000 152.640 ;
        RECT 4.400 150.640 56.000 152.000 ;
        RECT 4.400 150.600 55.600 150.640 ;
        RECT 3.990 149.960 55.600 150.600 ;
        RECT 4.400 149.240 55.600 149.960 ;
        RECT 4.400 148.560 56.000 149.240 ;
        RECT 3.990 147.240 56.000 148.560 ;
        RECT 4.400 146.560 56.000 147.240 ;
        RECT 4.400 145.840 55.600 146.560 ;
        RECT 3.990 145.200 55.600 145.840 ;
        RECT 4.400 145.160 55.600 145.200 ;
        RECT 4.400 143.800 56.000 145.160 ;
        RECT 3.990 143.160 56.000 143.800 ;
        RECT 4.400 141.760 55.600 143.160 ;
        RECT 3.990 141.120 56.000 141.760 ;
        RECT 4.400 139.720 56.000 141.120 ;
        RECT 3.990 139.080 56.000 139.720 ;
        RECT 4.400 137.680 55.600 139.080 ;
        RECT 3.990 137.040 56.000 137.680 ;
        RECT 4.400 135.680 56.000 137.040 ;
        RECT 4.400 135.640 55.600 135.680 ;
        RECT 3.990 135.000 55.600 135.640 ;
        RECT 4.400 134.280 55.600 135.000 ;
        RECT 4.400 133.600 56.000 134.280 ;
        RECT 3.990 132.280 56.000 133.600 ;
        RECT 4.400 131.600 56.000 132.280 ;
        RECT 4.400 130.880 55.600 131.600 ;
        RECT 3.990 130.240 55.600 130.880 ;
        RECT 4.400 130.200 55.600 130.240 ;
        RECT 4.400 128.840 56.000 130.200 ;
        RECT 3.990 128.200 56.000 128.840 ;
        RECT 4.400 127.520 56.000 128.200 ;
        RECT 4.400 126.800 55.600 127.520 ;
        RECT 3.990 126.160 55.600 126.800 ;
        RECT 4.400 126.120 55.600 126.160 ;
        RECT 4.400 124.760 56.000 126.120 ;
        RECT 3.990 124.120 56.000 124.760 ;
        RECT 4.400 122.720 55.600 124.120 ;
        RECT 3.990 122.080 56.000 122.720 ;
        RECT 4.400 120.680 56.000 122.080 ;
        RECT 3.990 120.040 56.000 120.680 ;
        RECT 3.990 119.360 55.600 120.040 ;
        RECT 4.400 118.640 55.600 119.360 ;
        RECT 4.400 117.960 56.000 118.640 ;
        RECT 3.990 117.320 56.000 117.960 ;
        RECT 4.400 116.640 56.000 117.320 ;
        RECT 4.400 115.920 55.600 116.640 ;
        RECT 3.990 115.280 55.600 115.920 ;
        RECT 4.400 115.240 55.600 115.280 ;
        RECT 4.400 113.880 56.000 115.240 ;
        RECT 3.990 113.240 56.000 113.880 ;
        RECT 4.400 112.560 56.000 113.240 ;
        RECT 4.400 111.840 55.600 112.560 ;
        RECT 3.990 111.200 55.600 111.840 ;
        RECT 4.400 111.160 55.600 111.200 ;
        RECT 4.400 109.800 56.000 111.160 ;
        RECT 3.990 109.160 56.000 109.800 ;
        RECT 4.400 108.480 56.000 109.160 ;
        RECT 4.400 107.760 55.600 108.480 ;
        RECT 3.990 107.080 55.600 107.760 ;
        RECT 3.990 106.440 56.000 107.080 ;
        RECT 4.400 105.080 56.000 106.440 ;
        RECT 4.400 105.040 55.600 105.080 ;
        RECT 3.990 104.400 55.600 105.040 ;
        RECT 4.400 103.680 55.600 104.400 ;
        RECT 4.400 103.000 56.000 103.680 ;
        RECT 3.990 102.360 56.000 103.000 ;
        RECT 4.400 101.000 56.000 102.360 ;
        RECT 4.400 100.960 55.600 101.000 ;
        RECT 3.990 100.320 55.600 100.960 ;
        RECT 4.400 99.600 55.600 100.320 ;
        RECT 4.400 98.920 56.000 99.600 ;
        RECT 3.990 98.280 56.000 98.920 ;
        RECT 4.400 97.600 56.000 98.280 ;
        RECT 4.400 96.880 55.600 97.600 ;
        RECT 3.990 96.240 55.600 96.880 ;
        RECT 4.400 96.200 55.600 96.240 ;
        RECT 4.400 94.840 56.000 96.200 ;
        RECT 3.990 93.520 56.000 94.840 ;
        RECT 4.400 92.120 55.600 93.520 ;
        RECT 3.990 91.480 56.000 92.120 ;
        RECT 4.400 90.080 56.000 91.480 ;
        RECT 3.990 89.440 56.000 90.080 ;
        RECT 4.400 88.040 55.600 89.440 ;
        RECT 3.990 87.400 56.000 88.040 ;
        RECT 4.400 86.040 56.000 87.400 ;
        RECT 4.400 86.000 55.600 86.040 ;
        RECT 3.990 85.360 55.600 86.000 ;
        RECT 4.400 84.640 55.600 85.360 ;
        RECT 4.400 83.960 56.000 84.640 ;
        RECT 3.990 83.320 56.000 83.960 ;
        RECT 4.400 81.960 56.000 83.320 ;
        RECT 4.400 81.920 55.600 81.960 ;
        RECT 3.990 80.600 55.600 81.920 ;
        RECT 4.400 80.560 55.600 80.600 ;
        RECT 4.400 79.200 56.000 80.560 ;
        RECT 3.990 78.560 56.000 79.200 ;
        RECT 4.400 77.160 55.600 78.560 ;
        RECT 3.990 76.520 56.000 77.160 ;
        RECT 4.400 75.120 56.000 76.520 ;
        RECT 3.990 74.480 56.000 75.120 ;
        RECT 4.400 73.080 55.600 74.480 ;
        RECT 3.990 72.440 56.000 73.080 ;
        RECT 4.400 71.040 56.000 72.440 ;
        RECT 3.990 70.400 56.000 71.040 ;
        RECT 4.400 69.000 55.600 70.400 ;
        RECT 3.990 68.360 56.000 69.000 ;
        RECT 4.400 67.000 56.000 68.360 ;
        RECT 4.400 66.960 55.600 67.000 ;
        RECT 3.990 65.640 55.600 66.960 ;
        RECT 4.400 65.600 55.600 65.640 ;
        RECT 4.400 64.240 56.000 65.600 ;
        RECT 3.990 63.600 56.000 64.240 ;
        RECT 4.400 62.920 56.000 63.600 ;
        RECT 4.400 62.200 55.600 62.920 ;
        RECT 3.990 61.560 55.600 62.200 ;
        RECT 4.400 61.520 55.600 61.560 ;
        RECT 4.400 60.160 56.000 61.520 ;
        RECT 3.990 59.520 56.000 60.160 ;
        RECT 4.400 58.120 55.600 59.520 ;
        RECT 3.990 57.480 56.000 58.120 ;
        RECT 4.400 56.080 56.000 57.480 ;
        RECT 3.990 55.440 56.000 56.080 ;
        RECT 4.400 54.040 55.600 55.440 ;
        RECT 3.990 52.720 56.000 54.040 ;
        RECT 4.400 51.360 56.000 52.720 ;
        RECT 4.400 51.320 55.600 51.360 ;
        RECT 3.990 50.680 55.600 51.320 ;
        RECT 4.400 49.960 55.600 50.680 ;
        RECT 4.400 49.280 56.000 49.960 ;
        RECT 3.990 48.640 56.000 49.280 ;
        RECT 4.400 47.960 56.000 48.640 ;
        RECT 4.400 47.240 55.600 47.960 ;
        RECT 3.990 46.600 55.600 47.240 ;
        RECT 4.400 46.560 55.600 46.600 ;
        RECT 4.400 45.200 56.000 46.560 ;
        RECT 3.990 44.560 56.000 45.200 ;
        RECT 4.400 43.880 56.000 44.560 ;
        RECT 4.400 43.160 55.600 43.880 ;
        RECT 3.990 42.520 55.600 43.160 ;
        RECT 4.400 42.480 55.600 42.520 ;
        RECT 4.400 41.120 56.000 42.480 ;
        RECT 3.990 40.480 56.000 41.120 ;
        RECT 3.990 39.800 55.600 40.480 ;
        RECT 4.400 39.080 55.600 39.800 ;
        RECT 4.400 38.400 56.000 39.080 ;
        RECT 3.990 37.760 56.000 38.400 ;
        RECT 4.400 36.400 56.000 37.760 ;
        RECT 4.400 36.360 55.600 36.400 ;
        RECT 3.990 35.720 55.600 36.360 ;
        RECT 4.400 35.000 55.600 35.720 ;
        RECT 4.400 34.320 56.000 35.000 ;
        RECT 3.990 33.680 56.000 34.320 ;
        RECT 4.400 32.320 56.000 33.680 ;
        RECT 4.400 32.280 55.600 32.320 ;
        RECT 3.990 31.640 55.600 32.280 ;
        RECT 4.400 30.920 55.600 31.640 ;
        RECT 4.400 30.240 56.000 30.920 ;
        RECT 3.990 29.600 56.000 30.240 ;
        RECT 4.400 28.920 56.000 29.600 ;
        RECT 4.400 28.200 55.600 28.920 ;
        RECT 3.990 27.520 55.600 28.200 ;
        RECT 3.990 26.880 56.000 27.520 ;
        RECT 4.400 25.480 56.000 26.880 ;
        RECT 3.990 24.840 56.000 25.480 ;
        RECT 4.400 23.440 55.600 24.840 ;
        RECT 3.990 22.800 56.000 23.440 ;
        RECT 4.400 21.440 56.000 22.800 ;
        RECT 4.400 21.400 55.600 21.440 ;
        RECT 3.990 20.760 55.600 21.400 ;
        RECT 4.400 20.040 55.600 20.760 ;
        RECT 4.400 19.360 56.000 20.040 ;
        RECT 3.990 18.720 56.000 19.360 ;
        RECT 4.400 17.360 56.000 18.720 ;
        RECT 4.400 17.320 55.600 17.360 ;
        RECT 3.990 16.680 55.600 17.320 ;
        RECT 4.400 15.960 55.600 16.680 ;
        RECT 4.400 15.280 56.000 15.960 ;
        RECT 3.990 13.960 56.000 15.280 ;
        RECT 4.400 13.280 56.000 13.960 ;
        RECT 4.400 12.560 55.600 13.280 ;
        RECT 3.990 11.920 55.600 12.560 ;
        RECT 4.400 11.880 55.600 11.920 ;
        RECT 4.400 10.520 56.000 11.880 ;
        RECT 3.990 9.880 56.000 10.520 ;
        RECT 4.400 8.480 55.600 9.880 ;
        RECT 3.990 7.840 56.000 8.480 ;
        RECT 4.400 6.440 56.000 7.840 ;
        RECT 3.990 5.800 56.000 6.440 ;
        RECT 4.400 4.400 55.600 5.800 ;
        RECT 3.990 3.760 56.000 4.400 ;
        RECT 4.400 2.400 56.000 3.760 ;
        RECT 4.400 2.360 55.600 2.400 ;
        RECT 3.990 1.720 55.600 2.360 ;
        RECT 4.400 1.000 55.600 1.720 ;
        RECT 4.400 0.855 56.000 1.000 ;
      LAYER met4 ;
        RECT 5.815 10.640 12.475 389.200 ;
        RECT 14.875 10.640 20.635 389.200 ;
        RECT 23.035 10.640 28.795 389.200 ;
        RECT 31.195 10.640 32.825 389.200 ;
  END
END wb_bridge_2way
END LIBRARY

