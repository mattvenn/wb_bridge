magic
tech sky130A
magscale 1 2
timestamp 1639997236
<< locali >>
rect 10977 76415 11011 77945
rect 949 74919 983 75905
rect 949 69343 983 74885
rect 11069 74537 11103 77333
rect 10977 74503 11103 74537
rect 3617 74103 3651 74409
rect 765 59755 799 66113
rect 857 61115 891 67881
rect 949 62339 983 67813
rect 857 59075 891 60809
rect 857 55675 891 59041
rect 949 55947 983 60673
rect 10977 55743 11011 74503
rect 11069 70567 11103 73525
rect 949 50167 983 51901
rect 10885 50167 10919 50405
rect 10977 50371 11011 54485
rect 6193 49623 6227 49793
rect 10977 48671 11011 50201
rect 11069 49351 11103 70397
rect 11161 69819 11195 72981
rect 11253 65551 11287 72165
rect 11345 70431 11379 74273
rect 11161 65517 11287 65551
rect 11161 49419 11195 65517
rect 11253 57511 11287 63937
rect 11069 49317 11195 49351
rect 10977 48637 11103 48671
rect 10977 45475 11011 48569
rect 11069 47039 11103 48637
rect 11069 45407 11103 46325
rect 10977 45373 11103 45407
rect 857 38811 891 44353
rect 949 41191 983 44217
rect 949 29699 983 34969
rect 3617 33983 3651 34153
rect 10977 31399 11011 45373
rect 11069 38539 11103 41565
rect 11161 40579 11195 49317
rect 11253 36771 11287 54145
rect 11345 37179 11379 64889
rect 11437 56763 11471 64481
rect 11529 55811 11563 61285
rect 11437 55777 11563 55811
rect 11437 34051 11471 55777
rect 11529 54111 11563 55709
rect 11621 54179 11655 62713
rect 11529 54077 11655 54111
rect 11529 50439 11563 53941
rect 11621 50439 11655 54077
rect 11713 53975 11747 56865
rect 11713 50371 11747 53669
rect 11529 50337 11747 50371
rect 11529 46359 11563 50337
rect 10977 29223 11011 30685
rect 11069 27387 11103 31297
rect 11161 27047 11195 31773
rect 11253 26503 11287 32385
rect 11529 31943 11563 46189
rect 11621 44523 11655 50269
rect 11713 49555 11747 50269
rect 11713 40375 11747 49385
rect 11805 41417 11839 69989
rect 11897 46223 11931 55641
rect 11805 41383 11931 41417
rect 11897 41191 11931 41383
rect 10977 16235 11011 19805
rect 10977 11339 11011 14365
rect 11069 12971 11103 17153
rect 11161 12903 11195 14977
rect 11069 12869 11195 12903
rect 11069 9163 11103 12869
rect 11253 12437 11287 16065
rect 11161 12403 11287 12437
rect 11161 8619 11195 12403
rect 11345 6917 11379 14297
rect 11161 6883 11379 6917
rect 11161 5219 11195 6883
<< viali >>
rect 10977 77945 11011 77979
rect 2697 77605 2731 77639
rect 9229 77605 9263 77639
rect 2513 77469 2547 77503
rect 3985 77469 4019 77503
rect 4629 77469 4663 77503
rect 5273 77469 5307 77503
rect 9413 77469 9447 77503
rect 10149 77469 10183 77503
rect 1777 77401 1811 77435
rect 1961 77401 1995 77435
rect 3801 77333 3835 77367
rect 4445 77333 4479 77367
rect 5089 77333 5123 77367
rect 9965 77333 9999 77367
rect 1409 76993 1443 77027
rect 2053 76993 2087 77027
rect 2697 76993 2731 77027
rect 3341 76993 3375 77027
rect 4169 76993 4203 77027
rect 10149 76993 10183 77027
rect 2881 76857 2915 76891
rect 1593 76789 1627 76823
rect 2237 76789 2271 76823
rect 3525 76789 3559 76823
rect 3985 76789 4019 76823
rect 9965 76789 9999 76823
rect 2237 76517 2271 76551
rect 1685 76381 1719 76415
rect 1869 76381 1903 76415
rect 2105 76381 2139 76415
rect 2973 76381 3007 76415
rect 10149 76381 10183 76415
rect 10977 76381 11011 76415
rect 11069 77333 11103 77367
rect 1961 76313 1995 76347
rect 2789 76245 2823 76279
rect 9965 76245 9999 76279
rect 1869 75973 1903 76007
rect 1961 75973 1995 76007
rect 949 75905 983 75939
rect 1685 75905 1719 75939
rect 2105 75905 2139 75939
rect 2973 75905 3007 75939
rect 10149 75905 10183 75939
rect 2237 75769 2271 75803
rect 2789 75701 2823 75735
rect 9965 75701 9999 75735
rect 2421 75429 2455 75463
rect 1409 75293 1443 75327
rect 2600 75293 2634 75327
rect 2697 75293 2731 75327
rect 2973 75293 3007 75327
rect 3985 75293 4019 75327
rect 10149 75293 10183 75327
rect 2789 75225 2823 75259
rect 1593 75157 1627 75191
rect 3801 75157 3835 75191
rect 9965 75157 9999 75191
rect 949 74885 983 74919
rect 3617 74885 3651 74919
rect 3709 74885 3743 74919
rect 1409 74817 1443 74851
rect 2600 74817 2634 74851
rect 2697 74817 2731 74851
rect 2789 74817 2823 74851
rect 2973 74817 3007 74851
rect 3433 74817 3467 74851
rect 3853 74817 3887 74851
rect 1593 74613 1627 74647
rect 2421 74613 2455 74647
rect 3985 74613 4019 74647
rect 3617 74409 3651 74443
rect 1961 74341 1995 74375
rect 2605 74341 2639 74375
rect 1409 74205 1443 74239
rect 1593 74205 1627 74239
rect 1685 74205 1719 74239
rect 1782 74205 1816 74239
rect 2743 74205 2777 74239
rect 2881 74205 2915 74239
rect 3157 74205 3191 74239
rect 2973 74137 3007 74171
rect 10149 74205 10183 74239
rect 3617 74069 3651 74103
rect 9965 74069 9999 74103
rect 1869 73797 1903 73831
rect 1633 73729 1667 73763
rect 1777 73729 1811 73763
rect 2053 73729 2087 73763
rect 2697 73729 2731 73763
rect 10149 73729 10183 73763
rect 1501 73593 1535 73627
rect 2513 73525 2547 73559
rect 9965 73525 9999 73559
rect 1409 73117 1443 73151
rect 2237 73117 2271 73151
rect 10149 73117 10183 73151
rect 1593 72981 1627 73015
rect 2053 72981 2087 73015
rect 9965 72981 9999 73015
rect 1409 72641 1443 72675
rect 1593 72437 1627 72471
rect 9965 72233 9999 72267
rect 1961 72165 1995 72199
rect 1409 72029 1443 72063
rect 1593 72029 1627 72063
rect 1829 72029 1863 72063
rect 10149 72029 10183 72063
rect 1685 71961 1719 71995
rect 9965 71689 9999 71723
rect 10149 71553 10183 71587
rect 1409 71485 1443 71519
rect 1685 71485 1719 71519
rect 1409 71009 1443 71043
rect 1685 70941 1719 70975
rect 2697 70941 2731 70975
rect 2881 70805 2915 70839
rect 9965 70601 9999 70635
rect 1685 70533 1719 70567
rect 2605 70533 2639 70567
rect 2461 70465 2495 70499
rect 2697 70465 2731 70499
rect 2881 70465 2915 70499
rect 3525 70465 3559 70499
rect 10149 70465 10183 70499
rect 2329 70329 2363 70363
rect 1593 70261 1627 70295
rect 3341 70261 3375 70295
rect 2421 69989 2455 70023
rect 1409 69853 1443 69887
rect 2600 69853 2634 69887
rect 2697 69853 2731 69887
rect 2973 69853 3007 69887
rect 3985 69853 4019 69887
rect 10149 69853 10183 69887
rect 2789 69785 2823 69819
rect 1593 69717 1627 69751
rect 3801 69717 3835 69751
rect 9965 69717 9999 69751
rect 1777 69445 1811 69479
rect 1639 69377 1673 69411
rect 1869 69377 1903 69411
rect 2053 69377 2087 69411
rect 3065 69377 3099 69411
rect 4261 69377 4295 69411
rect 10149 69377 10183 69411
rect 949 69309 983 69343
rect 2789 69309 2823 69343
rect 4077 69241 4111 69275
rect 1501 69173 1535 69207
rect 9965 69173 9999 69207
rect 2973 68833 3007 68867
rect 1409 68765 1443 68799
rect 3249 68765 3283 68799
rect 3985 68765 4019 68799
rect 1593 68629 1627 68663
rect 3801 68629 3835 68663
rect 3985 68425 4019 68459
rect 1961 68357 1995 68391
rect 2053 68357 2087 68391
rect 3065 68357 3099 68391
rect 3157 68357 3191 68391
rect 1777 68289 1811 68323
rect 2150 68289 2184 68323
rect 2881 68289 2915 68323
rect 3301 68289 3335 68323
rect 4169 68289 4203 68323
rect 10149 68289 10183 68323
rect 2329 68153 2363 68187
rect 9965 68153 9999 68187
rect 3433 68085 3467 68119
rect 857 67881 891 67915
rect 765 66113 799 66147
rect 949 67813 983 67847
rect 1409 67677 1443 67711
rect 1685 67677 1719 67711
rect 10149 67677 10183 67711
rect 2973 67609 3007 67643
rect 3157 67609 3191 67643
rect 9965 67541 9999 67575
rect 2973 67337 3007 67371
rect 2145 67269 2179 67303
rect 2001 67201 2035 67235
rect 2237 67201 2271 67235
rect 2421 67201 2455 67235
rect 3065 67201 3099 67235
rect 1869 67065 1903 67099
rect 1685 66589 1719 66623
rect 2329 66589 2363 66623
rect 2973 66589 3007 66623
rect 10149 66589 10183 66623
rect 1501 66453 1535 66487
rect 2145 66453 2179 66487
rect 2789 66453 2823 66487
rect 9965 66453 9999 66487
rect 1685 66113 1719 66147
rect 10149 66113 10183 66147
rect 1409 66045 1443 66079
rect 9965 65909 9999 65943
rect 1685 65501 1719 65535
rect 2145 65501 2179 65535
rect 2881 65501 2915 65535
rect 10149 65501 10183 65535
rect 1501 65365 1535 65399
rect 2329 65365 2363 65399
rect 3065 65365 3099 65399
rect 9965 65365 9999 65399
rect 1961 65093 1995 65127
rect 2053 65093 2087 65127
rect 1777 65025 1811 65059
rect 2150 65025 2184 65059
rect 3157 65025 3191 65059
rect 2881 64957 2915 64991
rect 2329 64889 2363 64923
rect 2605 64481 2639 64515
rect 9873 64481 9907 64515
rect 1685 64413 1719 64447
rect 2329 64413 2363 64447
rect 10149 64413 10183 64447
rect 1501 64277 1535 64311
rect 2237 64005 2271 64039
rect 2093 63937 2127 63971
rect 2329 63937 2363 63971
rect 2513 63937 2547 63971
rect 2973 63937 3007 63971
rect 3709 63937 3743 63971
rect 9873 63937 9907 63971
rect 10149 63869 10183 63903
rect 3893 63801 3927 63835
rect 1961 63733 1995 63767
rect 3157 63733 3191 63767
rect 1961 63529 1995 63563
rect 2605 63461 2639 63495
rect 1409 63325 1443 63359
rect 1829 63325 1863 63359
rect 2737 63325 2771 63359
rect 3019 63325 3053 63359
rect 3111 63325 3145 63359
rect 3801 63325 3835 63359
rect 1593 63257 1627 63291
rect 1685 63257 1719 63291
rect 2881 63257 2915 63291
rect 3985 63189 4019 63223
rect 9965 62985 9999 63019
rect 1685 62849 1719 62883
rect 2421 62849 2455 62883
rect 3157 62849 3191 62883
rect 4169 62849 4203 62883
rect 10149 62849 10183 62883
rect 2881 62781 2915 62815
rect 4261 62781 4295 62815
rect 1501 62645 1535 62679
rect 2237 62645 2271 62679
rect 1961 62441 1995 62475
rect 2605 62441 2639 62475
rect 949 62305 983 62339
rect 1409 62237 1443 62271
rect 1593 62237 1627 62271
rect 1685 62237 1719 62271
rect 1782 62237 1816 62271
rect 2737 62237 2771 62271
rect 3157 62237 3191 62271
rect 10149 62237 10183 62271
rect 2881 62169 2915 62203
rect 2973 62169 3007 62203
rect 9965 62101 9999 62135
rect 1978 61897 2012 61931
rect 1409 61761 1443 61795
rect 1593 61761 1627 61795
rect 1685 61761 1719 61795
rect 1782 61761 1816 61795
rect 2513 61761 2547 61795
rect 10149 61761 10183 61795
rect 2697 61557 2731 61591
rect 9965 61557 9999 61591
rect 1501 61285 1535 61319
rect 1680 61149 1714 61183
rect 1777 61149 1811 61183
rect 2053 61149 2087 61183
rect 2513 61149 2547 61183
rect 3801 61149 3835 61183
rect 857 61081 891 61115
rect 1869 61081 1903 61115
rect 2697 61013 2731 61047
rect 3985 61013 4019 61047
rect 765 59721 799 59755
rect 857 60809 891 60843
rect 2513 60741 2547 60775
rect 2605 60741 2639 60775
rect 857 59041 891 59075
rect 949 60673 983 60707
rect 1685 60673 1719 60707
rect 2329 60673 2363 60707
rect 2702 60673 2736 60707
rect 10149 60673 10183 60707
rect 9965 60537 9999 60571
rect 1501 60469 1535 60503
rect 2881 60469 2915 60503
rect 9965 60265 9999 60299
rect 2513 60129 2547 60163
rect 1685 60061 1719 60095
rect 2237 60061 2271 60095
rect 10149 60061 10183 60095
rect 1501 59925 1535 59959
rect 1685 59585 1719 59619
rect 2145 59585 2179 59619
rect 2329 59449 2363 59483
rect 1501 59381 1535 59415
rect 9965 59177 9999 59211
rect 2421 59041 2455 59075
rect 1685 58973 1719 59007
rect 2145 58973 2179 59007
rect 10149 58973 10183 59007
rect 1501 58837 1535 58871
rect 1685 58497 1719 58531
rect 10149 58497 10183 58531
rect 1501 58293 1535 58327
rect 9965 58293 9999 58327
rect 1961 58021 1995 58055
rect 1409 57885 1443 57919
rect 1829 57885 1863 57919
rect 2789 57885 2823 57919
rect 10149 57885 10183 57919
rect 1593 57817 1627 57851
rect 1685 57817 1719 57851
rect 2605 57749 2639 57783
rect 9965 57749 9999 57783
rect 2513 57545 2547 57579
rect 1593 57477 1627 57511
rect 2881 57477 2915 57511
rect 1409 57409 1443 57443
rect 1685 57409 1719 57443
rect 1829 57409 1863 57443
rect 2697 57409 2731 57443
rect 2789 57409 2823 57443
rect 3065 57409 3099 57443
rect 1961 57273 1995 57307
rect 9873 56865 9907 56899
rect 1685 56797 1719 56831
rect 2329 56797 2363 56831
rect 2697 56797 2731 56831
rect 10149 56797 10183 56831
rect 2513 56729 2547 56763
rect 2605 56729 2639 56763
rect 1501 56661 1535 56695
rect 2881 56661 2915 56695
rect 1501 56457 1535 56491
rect 2421 56389 2455 56423
rect 1685 56321 1719 56355
rect 2973 56321 3007 56355
rect 10149 56321 10183 56355
rect 2237 56185 2271 56219
rect 3157 56117 3191 56151
rect 9965 56117 9999 56151
rect 949 55913 983 55947
rect 3249 55845 3283 55879
rect 11345 74273 11379 74307
rect 11069 73525 11103 73559
rect 11069 70533 11103 70567
rect 11161 72981 11195 73015
rect 1685 55709 1719 55743
rect 2237 55709 2271 55743
rect 3801 55709 3835 55743
rect 10977 55709 11011 55743
rect 11069 70397 11103 70431
rect 857 55641 891 55675
rect 3065 55641 3099 55675
rect 1501 55573 1535 55607
rect 2421 55573 2455 55607
rect 3985 55573 4019 55607
rect 1685 55301 1719 55335
rect 1978 55301 2012 55335
rect 1409 55233 1443 55267
rect 1593 55233 1627 55267
rect 1829 55233 1863 55267
rect 2513 55233 2547 55267
rect 10149 55233 10183 55267
rect 2697 55097 2731 55131
rect 9965 55029 9999 55063
rect 1685 54621 1719 54655
rect 2421 54621 2455 54655
rect 10149 54621 10183 54655
rect 1501 54485 1535 54519
rect 2237 54485 2271 54519
rect 9965 54485 9999 54519
rect 10977 54485 11011 54519
rect 2973 54281 3007 54315
rect 1593 54145 1627 54179
rect 2881 54145 2915 54179
rect 3065 54145 3099 54179
rect 9873 54145 9907 54179
rect 1869 54077 1903 54111
rect 10057 53941 10091 53975
rect 1961 53669 1995 53703
rect 1409 53533 1443 53567
rect 1593 53533 1627 53567
rect 1829 53533 1863 53567
rect 2513 53533 2547 53567
rect 1685 53465 1719 53499
rect 2697 53397 2731 53431
rect 1685 53057 1719 53091
rect 2421 53057 2455 53091
rect 2881 53057 2915 53091
rect 9873 53057 9907 53091
rect 3065 52921 3099 52955
rect 1501 52853 1535 52887
rect 2237 52853 2271 52887
rect 10057 52853 10091 52887
rect 2145 52649 2179 52683
rect 2973 52649 3007 52683
rect 1685 52445 1719 52479
rect 2145 52445 2179 52479
rect 2329 52445 2363 52479
rect 2789 52445 2823 52479
rect 2973 52445 3007 52479
rect 9873 52445 9907 52479
rect 1501 52309 1535 52343
rect 10057 52309 10091 52343
rect 2973 52105 3007 52139
rect 3617 52105 3651 52139
rect 1685 51969 1719 52003
rect 2881 51969 2915 52003
rect 3077 51969 3111 52003
rect 3525 51969 3559 52003
rect 3709 51969 3743 52003
rect 949 51901 983 51935
rect 1501 51765 1535 51799
rect 2881 51561 2915 51595
rect 1685 51357 1719 51391
rect 2421 51357 2455 51391
rect 2881 51357 2915 51391
rect 3065 51357 3099 51391
rect 9873 51357 9907 51391
rect 1501 51221 1535 51255
rect 2237 51221 2271 51255
rect 10057 51221 10091 51255
rect 2237 51017 2271 51051
rect 2881 51017 2915 51051
rect 3525 50949 3559 50983
rect 1685 50881 1719 50915
rect 2145 50881 2179 50915
rect 2329 50881 2363 50915
rect 2789 50881 2823 50915
rect 2973 50881 3007 50915
rect 3433 50881 3467 50915
rect 3617 50881 3651 50915
rect 9873 50881 9907 50915
rect 1501 50677 1535 50711
rect 10057 50677 10091 50711
rect 3985 50473 4019 50507
rect 4629 50473 4663 50507
rect 1961 50405 1995 50439
rect 10885 50405 10919 50439
rect 2697 50337 2731 50371
rect 1409 50269 1443 50303
rect 1593 50269 1627 50303
rect 1777 50269 1811 50303
rect 2421 50269 2455 50303
rect 3801 50269 3835 50303
rect 3985 50269 4019 50303
rect 4445 50269 4479 50303
rect 4629 50269 4663 50303
rect 9873 50269 9907 50303
rect 1685 50201 1719 50235
rect 10977 50337 11011 50371
rect 949 50133 983 50167
rect 10057 50133 10091 50167
rect 10885 50133 10919 50167
rect 10977 50201 11011 50235
rect 1593 49861 1627 49895
rect 1685 49861 1719 49895
rect 1409 49793 1443 49827
rect 1777 49793 1811 49827
rect 2421 49793 2455 49827
rect 3341 49793 3375 49827
rect 3525 49793 3559 49827
rect 6193 49793 6227 49827
rect 3433 49725 3467 49759
rect 1961 49657 1995 49691
rect 2605 49589 2639 49623
rect 6193 49589 6227 49623
rect 1593 49181 1627 49215
rect 1685 49181 1719 49215
rect 1961 49181 1995 49215
rect 2697 49181 2731 49215
rect 3801 49181 3835 49215
rect 3985 49181 4019 49215
rect 9873 49181 9907 49215
rect 1777 49113 1811 49147
rect 1409 49045 1443 49079
rect 2513 49045 2547 49079
rect 3893 49045 3927 49079
rect 10057 49045 10091 49079
rect 2237 48841 2271 48875
rect 1685 48705 1719 48739
rect 2421 48705 2455 48739
rect 3249 48705 3283 48739
rect 3433 48705 3467 48739
rect 9873 48705 9907 48739
rect 11161 69785 11195 69819
rect 11253 72165 11287 72199
rect 11345 70397 11379 70431
rect 11805 69989 11839 70023
rect 11345 64889 11379 64923
rect 11253 63937 11287 63971
rect 11253 57477 11287 57511
rect 11161 49385 11195 49419
rect 11253 54145 11287 54179
rect 3341 48637 3375 48671
rect 10977 48569 11011 48603
rect 1501 48501 1535 48535
rect 10057 48501 10091 48535
rect 2973 48229 3007 48263
rect 2237 48161 2271 48195
rect 1685 48093 1719 48127
rect 2145 48093 2179 48127
rect 2329 48093 2363 48127
rect 2789 48093 2823 48127
rect 2973 48093 3007 48127
rect 1501 47957 1535 47991
rect 2881 47753 2915 47787
rect 1685 47617 1719 47651
rect 2421 47617 2455 47651
rect 3065 47617 3099 47651
rect 9873 47617 9907 47651
rect 10057 47481 10091 47515
rect 1501 47413 1535 47447
rect 2237 47413 2271 47447
rect 2145 47209 2179 47243
rect 2973 47209 3007 47243
rect 1685 47005 1719 47039
rect 2145 47005 2179 47039
rect 2329 47005 2363 47039
rect 2973 47005 3007 47039
rect 9873 47005 9907 47039
rect 1501 46869 1535 46903
rect 10057 46869 10091 46903
rect 2329 46665 2363 46699
rect 2973 46665 3007 46699
rect 1685 46529 1719 46563
rect 2237 46529 2271 46563
rect 2421 46529 2455 46563
rect 2881 46529 2915 46563
rect 3065 46529 3099 46563
rect 9873 46529 9907 46563
rect 1501 46325 1535 46359
rect 10057 46325 10091 46359
rect 1685 45985 1719 46019
rect 1777 45917 1811 45951
rect 2053 45917 2087 45951
rect 2513 45917 2547 45951
rect 2697 45781 2731 45815
rect 11069 47005 11103 47039
rect 1685 45441 1719 45475
rect 9873 45441 9907 45475
rect 10977 45441 11011 45475
rect 11069 46325 11103 46359
rect 3433 45373 3467 45407
rect 3709 45373 3743 45407
rect 1501 45237 1535 45271
rect 10057 45237 10091 45271
rect 1501 44897 1535 44931
rect 1685 44829 1719 44863
rect 1869 44829 1903 44863
rect 2605 44829 2639 44863
rect 3065 44829 3099 44863
rect 3249 44829 3283 44863
rect 3801 44829 3835 44863
rect 3985 44829 4019 44863
rect 9873 44829 9907 44863
rect 3157 44761 3191 44795
rect 2421 44693 2455 44727
rect 3893 44693 3927 44727
rect 10057 44693 10091 44727
rect 3157 44489 3191 44523
rect 3801 44489 3835 44523
rect 4445 44489 4479 44523
rect 857 44353 891 44387
rect 1501 44353 1535 44387
rect 1685 44353 1719 44387
rect 2329 44353 2363 44387
rect 3065 44353 3099 44387
rect 3249 44353 3283 44387
rect 3709 44353 3743 44387
rect 3893 44353 3927 44387
rect 4353 44353 4387 44387
rect 4537 44353 4571 44387
rect 949 44217 983 44251
rect 1777 44217 1811 44251
rect 2513 44149 2547 44183
rect 1593 43945 1627 43979
rect 4445 43877 4479 43911
rect 1409 43741 1443 43775
rect 2421 43741 2455 43775
rect 2881 43741 2915 43775
rect 4261 43741 4295 43775
rect 4905 43741 4939 43775
rect 5089 43741 5123 43775
rect 9873 43741 9907 43775
rect 2237 43605 2271 43639
rect 3065 43605 3099 43639
rect 4997 43605 5031 43639
rect 10057 43605 10091 43639
rect 2237 43401 2271 43435
rect 1685 43265 1719 43299
rect 2145 43265 2179 43299
rect 2329 43265 2363 43299
rect 3065 43265 3099 43299
rect 9873 43265 9907 43299
rect 2789 43197 2823 43231
rect 1501 43061 1535 43095
rect 10057 43061 10091 43095
rect 1685 42653 1719 42687
rect 2421 42653 2455 42687
rect 9873 42653 9907 42687
rect 1501 42517 1535 42551
rect 2237 42517 2271 42551
rect 10057 42517 10091 42551
rect 3433 42245 3467 42279
rect 4169 42245 4203 42279
rect 4353 42245 4387 42279
rect 1685 42177 1719 42211
rect 3617 42041 3651 42075
rect 1501 41973 1535 42007
rect 2145 41769 2179 41803
rect 4077 41769 4111 41803
rect 1685 41565 1719 41599
rect 2329 41565 2363 41599
rect 3893 41565 3927 41599
rect 4077 41565 4111 41599
rect 9873 41565 9907 41599
rect 1501 41429 1535 41463
rect 10057 41429 10091 41463
rect 1777 41225 1811 41259
rect 949 41157 983 41191
rect 1501 41089 1535 41123
rect 1777 41089 1811 41123
rect 2605 41089 2639 41123
rect 9873 41089 9907 41123
rect 2421 40953 2455 40987
rect 10057 40885 10091 40919
rect 3801 40681 3835 40715
rect 1685 40477 1719 40511
rect 2145 40477 2179 40511
rect 2881 40477 2915 40511
rect 3801 40477 3835 40511
rect 3985 40477 4019 40511
rect 1501 40341 1535 40375
rect 2329 40341 2363 40375
rect 3065 40341 3099 40375
rect 1961 40137 1995 40171
rect 2789 40069 2823 40103
rect 1961 40001 1995 40035
rect 2237 40001 2271 40035
rect 2973 40001 3007 40035
rect 3433 40001 3467 40035
rect 3617 40001 3651 40035
rect 4083 40001 4117 40035
rect 4261 40001 4295 40035
rect 9873 40001 9907 40035
rect 4169 39933 4203 39967
rect 3433 39865 3467 39899
rect 10057 39865 10091 39899
rect 3801 39593 3835 39627
rect 4537 39457 4571 39491
rect 1685 39389 1719 39423
rect 2421 39389 2455 39423
rect 3157 39389 3191 39423
rect 3801 39389 3835 39423
rect 3985 39389 4019 39423
rect 4445 39389 4479 39423
rect 4629 39389 4663 39423
rect 9873 39389 9907 39423
rect 1501 39253 1535 39287
rect 2237 39253 2271 39287
rect 2973 39253 3007 39287
rect 10057 39253 10091 39287
rect 4353 39049 4387 39083
rect 1685 38981 1719 39015
rect 1869 38913 1903 38947
rect 2053 38913 2087 38947
rect 2973 38913 3007 38947
rect 3617 38913 3651 38947
rect 3801 38913 3835 38947
rect 4261 38913 4295 38947
rect 4445 38913 4479 38947
rect 9873 38913 9907 38947
rect 3709 38845 3743 38879
rect 857 38777 891 38811
rect 3157 38777 3191 38811
rect 10057 38709 10091 38743
rect 2881 38505 2915 38539
rect 3985 38505 4019 38539
rect 2237 38301 2271 38335
rect 3801 38301 3835 38335
rect 3985 38301 4019 38335
rect 2973 38233 3007 38267
rect 2145 38165 2179 38199
rect 2329 37961 2363 37995
rect 1685 37825 1719 37859
rect 2513 37825 2547 37859
rect 9873 37825 9907 37859
rect 1501 37621 1535 37655
rect 10057 37621 10091 37655
rect 2329 37417 2363 37451
rect 1501 37213 1535 37247
rect 1685 37213 1719 37247
rect 2513 37213 2547 37247
rect 2973 37213 3007 37247
rect 3065 37213 3099 37247
rect 9873 37213 9907 37247
rect 1685 37077 1719 37111
rect 10057 37077 10091 37111
rect 3709 36873 3743 36907
rect 1685 36737 1719 36771
rect 2421 36737 2455 36771
rect 2881 36737 2915 36771
rect 3617 36737 3651 36771
rect 3801 36737 3835 36771
rect 3065 36601 3099 36635
rect 1501 36533 1535 36567
rect 2237 36533 2271 36567
rect 3985 36329 4019 36363
rect 1685 36125 1719 36159
rect 3801 36125 3835 36159
rect 3985 36125 4019 36159
rect 9873 36125 9907 36159
rect 1501 35989 1535 36023
rect 10057 35989 10091 36023
rect 1777 35785 1811 35819
rect 1593 35649 1627 35683
rect 1777 35649 1811 35683
rect 2513 35649 2547 35683
rect 2789 35649 2823 35683
rect 3433 35649 3467 35683
rect 9873 35649 9907 35683
rect 3709 35581 3743 35615
rect 2513 35513 2547 35547
rect 10057 35445 10091 35479
rect 3249 35241 3283 35275
rect 2513 35173 2547 35207
rect 1685 35037 1719 35071
rect 2237 35037 2271 35071
rect 2421 35037 2455 35071
rect 3065 35037 3099 35071
rect 3249 35037 3283 35071
rect 9873 35037 9907 35071
rect 949 34969 983 35003
rect 1501 34901 1535 34935
rect 10057 34901 10091 34935
rect 1501 34697 1535 34731
rect 2605 34629 2639 34663
rect 1593 34561 1627 34595
rect 2237 34561 2271 34595
rect 2421 34561 2455 34595
rect 3065 34561 3099 34595
rect 3249 34357 3283 34391
rect 3617 34153 3651 34187
rect 3985 34153 4019 34187
rect 3065 34085 3099 34119
rect 1685 33949 1719 33983
rect 2145 33949 2179 33983
rect 2881 33949 2915 33983
rect 3617 33949 3651 33983
rect 3801 33949 3835 33983
rect 3985 33949 4019 33983
rect 9873 33949 9907 33983
rect 1501 33813 1535 33847
rect 2329 33813 2363 33847
rect 10057 33813 10091 33847
rect 2513 33609 2547 33643
rect 3157 33609 3191 33643
rect 1685 33473 1719 33507
rect 2329 33473 2363 33507
rect 2605 33473 2639 33507
rect 3065 33473 3099 33507
rect 3249 33473 3283 33507
rect 9873 33473 9907 33507
rect 1501 33269 1535 33303
rect 10057 33269 10091 33303
rect 2881 33065 2915 33099
rect 3801 33065 3835 33099
rect 1685 32861 1719 32895
rect 2145 32861 2179 32895
rect 2881 32861 2915 32895
rect 3065 32861 3099 32895
rect 3801 32861 3835 32895
rect 3985 32861 4019 32895
rect 1501 32725 1535 32759
rect 2329 32725 2363 32759
rect 1501 32521 1535 32555
rect 3341 32521 3375 32555
rect 2421 32453 2455 32487
rect 1409 32385 1443 32419
rect 1593 32385 1627 32419
rect 2145 32385 2179 32419
rect 2237 32385 2271 32419
rect 3249 32385 3283 32419
rect 3433 32385 3467 32419
rect 9873 32385 9907 32419
rect 10057 32249 10091 32283
rect 1593 31977 1627 32011
rect 3985 31977 4019 32011
rect 1777 31773 1811 31807
rect 2237 31773 2271 31807
rect 3801 31773 3835 31807
rect 3985 31773 4019 31807
rect 9873 31773 9907 31807
rect 2421 31637 2455 31671
rect 10057 31637 10091 31671
rect 11069 41565 11103 41599
rect 11161 40545 11195 40579
rect 11069 38505 11103 38539
rect 11437 64481 11471 64515
rect 11621 62713 11655 62747
rect 11437 56729 11471 56763
rect 11529 61285 11563 61319
rect 11345 37145 11379 37179
rect 11253 36737 11287 36771
rect 11529 55709 11563 55743
rect 11621 54145 11655 54179
rect 11713 56865 11747 56899
rect 11529 53941 11563 53975
rect 11529 50405 11563 50439
rect 11713 53941 11747 53975
rect 11621 50405 11655 50439
rect 11713 53669 11747 53703
rect 11529 46325 11563 46359
rect 11621 50269 11655 50303
rect 11437 34017 11471 34051
rect 11529 46189 11563 46223
rect 11253 32385 11287 32419
rect 1501 31365 1535 31399
rect 10977 31365 11011 31399
rect 11161 31773 11195 31807
rect 1777 31297 1811 31331
rect 2237 31297 2271 31331
rect 9873 31297 9907 31331
rect 11069 31297 11103 31331
rect 2421 31093 2455 31127
rect 10057 31093 10091 31127
rect 1685 30685 1719 30719
rect 2329 30685 2363 30719
rect 10149 30685 10183 30719
rect 10977 30685 11011 30719
rect 1501 30549 1535 30583
rect 2145 30549 2179 30583
rect 1593 30277 1627 30311
rect 1685 30209 1719 30243
rect 2145 30209 2179 30243
rect 2973 30209 3007 30243
rect 9873 30209 9907 30243
rect 2329 30073 2363 30107
rect 2789 30005 2823 30039
rect 10057 30005 10091 30039
rect 1593 29801 1627 29835
rect 2237 29801 2271 29835
rect 2881 29801 2915 29835
rect 949 29665 983 29699
rect 1777 29597 1811 29631
rect 2421 29597 2455 29631
rect 3065 29597 3099 29631
rect 3617 29257 3651 29291
rect 10977 29189 11011 29223
rect 2053 29121 2087 29155
rect 2237 29121 2271 29155
rect 2881 29121 2915 29155
rect 3065 29121 3099 29155
rect 3801 29121 3835 29155
rect 2329 29053 2363 29087
rect 2881 28985 2915 29019
rect 10149 28917 10183 28951
rect 2605 28713 2639 28747
rect 2053 28645 2087 28679
rect 2053 28509 2087 28543
rect 2789 28509 2823 28543
rect 3985 28509 4019 28543
rect 3801 28373 3835 28407
rect 3801 28169 3835 28203
rect 1501 28101 1535 28135
rect 1777 28033 1811 28067
rect 2329 28033 2363 28067
rect 2513 28033 2547 28067
rect 3341 28033 3375 28067
rect 3985 28033 4019 28067
rect 2329 27897 2363 27931
rect 3157 27829 3191 27863
rect 2329 27557 2363 27591
rect 3985 27557 4019 27591
rect 3157 27489 3191 27523
rect 10149 27489 10183 27523
rect 1409 27421 1443 27455
rect 2145 27421 2179 27455
rect 2329 27421 2363 27455
rect 3065 27421 3099 27455
rect 3249 27421 3283 27455
rect 3807 27421 3841 27455
rect 3985 27421 4019 27455
rect 11069 27353 11103 27387
rect 1593 27285 1627 27319
rect 4537 27081 4571 27115
rect 1593 27013 1627 27047
rect 3157 27013 3191 27047
rect 3985 27013 4019 27047
rect 11161 27013 11195 27047
rect 1869 26945 1903 26979
rect 2513 26945 2547 26979
rect 2605 26945 2639 26979
rect 3341 26945 3375 26979
rect 3893 26945 3927 26979
rect 4077 26945 4111 26979
rect 4721 26945 4755 26979
rect 10149 26945 10183 26979
rect 2421 26809 2455 26843
rect 3801 26537 3835 26571
rect 11713 50269 11747 50303
rect 11713 49521 11747 49555
rect 11621 44489 11655 44523
rect 11713 49385 11747 49419
rect 11897 55641 11931 55675
rect 11897 46189 11931 46223
rect 11897 41157 11931 41191
rect 11713 40341 11747 40375
rect 11529 31909 11563 31943
rect 3157 26469 3191 26503
rect 11253 26469 11287 26503
rect 1409 26333 1443 26367
rect 2053 26333 2087 26367
rect 2973 26333 3007 26367
rect 3157 26333 3191 26367
rect 3985 26333 4019 26367
rect 1593 26197 1627 26231
rect 2237 26197 2271 26231
rect 2145 25925 2179 25959
rect 1869 25857 1903 25891
rect 2789 25857 2823 25891
rect 2605 25653 2639 25687
rect 2329 25449 2363 25483
rect 10149 25449 10183 25483
rect 1869 25381 1903 25415
rect 1869 25245 1903 25279
rect 2329 25245 2363 25279
rect 3249 25245 3283 25279
rect 3065 25109 3099 25143
rect 3065 24837 3099 24871
rect 1409 24769 1443 24803
rect 2329 24769 2363 24803
rect 3433 24769 3467 24803
rect 10149 24769 10183 24803
rect 1593 24633 1627 24667
rect 2329 24565 2363 24599
rect 2421 24361 2455 24395
rect 10149 24361 10183 24395
rect 1409 24157 1443 24191
rect 2237 24157 2271 24191
rect 3157 24157 3191 24191
rect 1593 24021 1627 24055
rect 2973 24021 3007 24055
rect 2237 23749 2271 23783
rect 1409 23681 1443 23715
rect 2513 23681 2547 23715
rect 9873 23681 9907 23715
rect 1593 23477 1627 23511
rect 10057 23477 10091 23511
rect 1593 23273 1627 23307
rect 3065 23273 3099 23307
rect 9505 23273 9539 23307
rect 10149 23273 10183 23307
rect 2329 23205 2363 23239
rect 1593 23069 1627 23103
rect 2145 23069 2179 23103
rect 2973 23069 3007 23103
rect 9321 23069 9355 23103
rect 2421 22729 2455 22763
rect 1869 22593 1903 22627
rect 2513 22593 2547 22627
rect 3157 22593 3191 22627
rect 9873 22593 9907 22627
rect 2973 22457 3007 22491
rect 1869 22389 1903 22423
rect 10057 22389 10091 22423
rect 3801 22185 3835 22219
rect 1961 22049 1995 22083
rect 2237 21981 2271 22015
rect 2881 21981 2915 22015
rect 3985 21981 4019 22015
rect 9873 21981 9907 22015
rect 2697 21845 2731 21879
rect 10057 21845 10091 21879
rect 1869 21641 1903 21675
rect 3249 21573 3283 21607
rect 1961 21505 1995 21539
rect 2881 21505 2915 21539
rect 3893 21505 3927 21539
rect 2513 21369 2547 21403
rect 3709 21301 3743 21335
rect 1961 21097 1995 21131
rect 3801 21097 3835 21131
rect 2881 21029 2915 21063
rect 2053 20893 2087 20927
rect 3985 20893 4019 20927
rect 9873 20893 9907 20927
rect 2513 20825 2547 20859
rect 2697 20825 2731 20859
rect 10057 20757 10091 20791
rect 1593 20553 1627 20587
rect 2605 20553 2639 20587
rect 3893 20553 3927 20587
rect 9413 20553 9447 20587
rect 1685 20417 1719 20451
rect 2789 20417 2823 20451
rect 3433 20417 3467 20451
rect 4077 20417 4111 20451
rect 9229 20417 9263 20451
rect 9873 20417 9907 20451
rect 3249 20213 3283 20247
rect 10057 20213 10091 20247
rect 1961 20009 1995 20043
rect 2605 20009 2639 20043
rect 2053 19805 2087 19839
rect 2697 19805 2731 19839
rect 9873 19805 9907 19839
rect 10977 19805 11011 19839
rect 4353 19737 4387 19771
rect 4261 19669 4295 19703
rect 10057 19669 10091 19703
rect 2329 19465 2363 19499
rect 2881 19465 2915 19499
rect 9965 19465 9999 19499
rect 1409 19329 1443 19363
rect 2421 19329 2455 19363
rect 3065 19329 3099 19363
rect 10149 19329 10183 19363
rect 1593 19125 1627 19159
rect 1869 18921 1903 18955
rect 9413 18921 9447 18955
rect 3065 18853 3099 18887
rect 1961 18717 1995 18751
rect 2605 18717 2639 18751
rect 3249 18717 3283 18751
rect 9229 18717 9263 18751
rect 9873 18717 9907 18751
rect 2421 18581 2455 18615
rect 10057 18581 10091 18615
rect 2145 18377 2179 18411
rect 2697 18377 2731 18411
rect 1593 18241 1627 18275
rect 2237 18241 2271 18275
rect 2881 18241 2915 18275
rect 9873 18241 9907 18275
rect 1501 18173 1535 18207
rect 10057 18037 10091 18071
rect 1777 17833 1811 17867
rect 9873 17833 9907 17867
rect 2881 17697 2915 17731
rect 1685 17629 1719 17663
rect 2513 17629 2547 17663
rect 10057 17629 10091 17663
rect 2605 17493 2639 17527
rect 2697 17493 2731 17527
rect 2881 17493 2915 17527
rect 2697 17289 2731 17323
rect 1409 17153 1443 17187
rect 2237 17153 2271 17187
rect 2881 17153 2915 17187
rect 9873 17153 9907 17187
rect 10057 17017 10091 17051
rect 1593 16949 1627 16983
rect 2053 16949 2087 16983
rect 3065 16745 3099 16779
rect 2973 16609 3007 16643
rect 1409 16541 1443 16575
rect 2789 16541 2823 16575
rect 9229 16541 9263 16575
rect 9873 16541 9907 16575
rect 3065 16473 3099 16507
rect 1593 16405 1627 16439
rect 2605 16405 2639 16439
rect 9413 16405 9447 16439
rect 10057 16405 10091 16439
rect 1961 16201 1995 16235
rect 9413 16201 9447 16235
rect 10977 16201 11011 16235
rect 11069 17153 11103 17187
rect 1501 16065 1535 16099
rect 1777 16065 1811 16099
rect 2605 16065 2639 16099
rect 3249 16065 3283 16099
rect 9229 16065 9263 16099
rect 9873 16065 9907 16099
rect 1685 15997 1719 16031
rect 3065 15929 3099 15963
rect 1777 15861 1811 15895
rect 2421 15861 2455 15895
rect 10057 15861 10091 15895
rect 1501 15657 1535 15691
rect 2697 15657 2731 15691
rect 9965 15657 9999 15691
rect 2789 15521 2823 15555
rect 1409 15453 1443 15487
rect 1593 15453 1627 15487
rect 2414 15453 2448 15487
rect 10149 15453 10183 15487
rect 2513 15317 2547 15351
rect 2605 15317 2639 15351
rect 1409 15113 1443 15147
rect 2605 15113 2639 15147
rect 9413 15113 9447 15147
rect 3525 15045 3559 15079
rect 1593 14977 1627 15011
rect 1869 14977 1903 15011
rect 2421 14977 2455 15011
rect 2697 14977 2731 15011
rect 3157 14977 3191 15011
rect 3341 14977 3375 15011
rect 9229 14977 9263 15011
rect 9873 14977 9907 15011
rect 1685 14909 1719 14943
rect 1869 14773 1903 14807
rect 10057 14773 10091 14807
rect 4445 14569 4479 14603
rect 3801 14501 3835 14535
rect 2145 14365 2179 14399
rect 2329 14365 2363 14399
rect 3065 14365 3099 14399
rect 3249 14365 3283 14399
rect 3985 14365 4019 14399
rect 4629 14365 4663 14399
rect 9873 14365 9907 14399
rect 10977 14365 11011 14399
rect 3157 14297 3191 14331
rect 2237 14229 2271 14263
rect 10057 14229 10091 14263
rect 2605 14025 2639 14059
rect 3341 14025 3375 14059
rect 3985 14025 4019 14059
rect 2053 13957 2087 13991
rect 1869 13889 1903 13923
rect 2513 13889 2547 13923
rect 3157 13889 3191 13923
rect 3801 13889 3835 13923
rect 4629 13889 4663 13923
rect 4445 13753 4479 13787
rect 2881 13481 2915 13515
rect 1685 13345 1719 13379
rect 1409 13277 1443 13311
rect 2789 13277 2823 13311
rect 2973 13277 3007 13311
rect 4353 13277 4387 13311
rect 9873 13277 9907 13311
rect 4169 13209 4203 13243
rect 10057 13141 10091 13175
rect 9413 12937 9447 12971
rect 1685 12801 1719 12835
rect 9229 12801 9263 12835
rect 9873 12801 9907 12835
rect 1409 12733 1443 12767
rect 2697 12733 2731 12767
rect 2973 12733 3007 12767
rect 10057 12597 10091 12631
rect 2789 12393 2823 12427
rect 1685 12257 1719 12291
rect 1409 12189 1443 12223
rect 2973 12189 3007 12223
rect 9873 12189 9907 12223
rect 10057 12053 10091 12087
rect 2789 11849 2823 11883
rect 9965 11849 9999 11883
rect 1685 11713 1719 11747
rect 2973 11713 3007 11747
rect 10149 11713 10183 11747
rect 1409 11645 1443 11679
rect 11253 16065 11287 16099
rect 11069 12937 11103 12971
rect 11161 14977 11195 15011
rect 2789 11305 2823 11339
rect 9413 11305 9447 11339
rect 10977 11305 11011 11339
rect 1685 11169 1719 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 3801 11101 3835 11135
rect 9229 11101 9263 11135
rect 9873 11101 9907 11135
rect 3985 10965 4019 10999
rect 10057 10965 10091 10999
rect 1685 10625 1719 10659
rect 2697 10625 2731 10659
rect 9873 10625 9907 10659
rect 1409 10557 1443 10591
rect 2881 10421 2915 10455
rect 10057 10421 10091 10455
rect 2789 10217 2823 10251
rect 1685 10081 1719 10115
rect 1409 10013 1443 10047
rect 2973 10013 3007 10047
rect 2789 9673 2823 9707
rect 2697 9537 2731 9571
rect 2911 9537 2945 9571
rect 9873 9537 9907 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3065 9469 3099 9503
rect 2973 9401 3007 9435
rect 10057 9401 10091 9435
rect 1593 9129 1627 9163
rect 9413 9129 9447 9163
rect 11069 9129 11103 9163
rect 11345 14297 11379 14331
rect 2421 9061 2455 9095
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 2881 8925 2915 8959
rect 3801 8925 3835 8959
rect 9229 8925 9263 8959
rect 9873 8925 9907 8959
rect 3065 8789 3099 8823
rect 3985 8789 4019 8823
rect 10057 8789 10091 8823
rect 1593 8585 1627 8619
rect 9413 8585 9447 8619
rect 11161 8585 11195 8619
rect 1409 8449 1443 8483
rect 2513 8449 2547 8483
rect 9229 8449 9263 8483
rect 9873 8449 9907 8483
rect 2697 8313 2731 8347
rect 10057 8245 10091 8279
rect 1685 7905 1719 7939
rect 1409 7837 1443 7871
rect 3065 7837 3099 7871
rect 3249 7837 3283 7871
rect 3157 7701 3191 7735
rect 2881 7497 2915 7531
rect 1409 7361 1443 7395
rect 2697 7361 2731 7395
rect 3433 7361 3467 7395
rect 3617 7361 3651 7395
rect 9873 7361 9907 7395
rect 1685 7293 1719 7327
rect 3617 7157 3651 7191
rect 10057 7157 10091 7191
rect 2145 6817 2179 6851
rect 2973 6749 3007 6783
rect 3801 6749 3835 6783
rect 9873 6749 9907 6783
rect 1869 6681 1903 6715
rect 2789 6613 2823 6647
rect 3985 6613 4019 6647
rect 10057 6613 10091 6647
rect 3249 6409 3283 6443
rect 1961 6273 1995 6307
rect 2605 6273 2639 6307
rect 3433 6273 3467 6307
rect 2789 6137 2823 6171
rect 2145 6069 2179 6103
rect 2789 5865 2823 5899
rect 3801 5865 3835 5899
rect 1501 5797 1535 5831
rect 1685 5661 1719 5695
rect 2145 5661 2179 5695
rect 2973 5661 3007 5695
rect 3985 5661 4019 5695
rect 9873 5661 9907 5695
rect 2329 5525 2363 5559
rect 10057 5525 10091 5559
rect 1961 5321 1995 5355
rect 2053 5185 2087 5219
rect 2973 5185 3007 5219
rect 3157 5185 3191 5219
rect 9873 5185 9907 5219
rect 11161 5185 11195 5219
rect 3157 4981 3191 5015
rect 10057 4981 10091 5015
rect 3801 4777 3835 4811
rect 1593 4709 1627 4743
rect 1409 4573 1443 4607
rect 2421 4573 2455 4607
rect 3065 4573 3099 4607
rect 3985 4573 4019 4607
rect 9873 4573 9907 4607
rect 2605 4437 2639 4471
rect 3249 4437 3283 4471
rect 10057 4437 10091 4471
rect 1869 4097 1903 4131
rect 2145 4097 2179 4131
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 3341 4097 3375 4131
rect 3525 4097 3559 4131
rect 4169 4097 4203 4131
rect 3525 3961 3559 3995
rect 3985 3893 4019 3927
rect 2237 3689 2271 3723
rect 1501 3621 1535 3655
rect 1685 3485 1719 3519
rect 2329 3485 2363 3519
rect 2973 3485 3007 3519
rect 3157 3485 3191 3519
rect 9873 3485 9907 3519
rect 3065 3349 3099 3383
rect 10057 3349 10091 3383
rect 3985 3145 4019 3179
rect 1685 3009 1719 3043
rect 2881 3009 2915 3043
rect 3525 3009 3559 3043
rect 4169 3009 4203 3043
rect 9137 3009 9171 3043
rect 9873 3009 9907 3043
rect 1409 2941 1443 2975
rect 2697 2873 2731 2907
rect 3341 2873 3375 2907
rect 9321 2805 9355 2839
rect 10057 2805 10091 2839
rect 1593 2601 1627 2635
rect 2237 2601 2271 2635
rect 2697 2601 2731 2635
rect 3801 2601 3835 2635
rect 4445 2601 4479 2635
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 2881 2397 2915 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 9137 2397 9171 2431
rect 9873 2397 9907 2431
rect 9321 2261 9355 2295
rect 10057 2261 10091 2295
<< metal1 >>
rect 10962 77976 10968 77988
rect 10923 77948 10968 77976
rect 10962 77936 10968 77948
rect 11020 77936 11026 77988
rect 1104 77818 10856 77840
rect 1104 77766 2582 77818
rect 2634 77766 2646 77818
rect 2698 77766 2710 77818
rect 2762 77766 2774 77818
rect 2826 77766 2838 77818
rect 2890 77766 5845 77818
rect 5897 77766 5909 77818
rect 5961 77766 5973 77818
rect 6025 77766 6037 77818
rect 6089 77766 6101 77818
rect 6153 77766 9109 77818
rect 9161 77766 9173 77818
rect 9225 77766 9237 77818
rect 9289 77766 9301 77818
rect 9353 77766 9365 77818
rect 9417 77766 10856 77818
rect 1104 77744 10856 77766
rect 2685 77639 2743 77645
rect 2685 77605 2697 77639
rect 2731 77636 2743 77639
rect 3234 77636 3240 77648
rect 2731 77608 3240 77636
rect 2731 77605 2743 77608
rect 2685 77599 2743 77605
rect 3234 77596 3240 77608
rect 3292 77596 3298 77648
rect 4706 77596 4712 77648
rect 4764 77636 4770 77648
rect 9217 77639 9275 77645
rect 9217 77636 9229 77639
rect 4764 77608 9229 77636
rect 4764 77596 4770 77608
rect 9217 77605 9229 77608
rect 9263 77605 9275 77639
rect 9217 77599 9275 77605
rect 3050 77528 3056 77580
rect 3108 77568 3114 77580
rect 3108 77540 5304 77568
rect 3108 77528 3114 77540
rect 2498 77500 2504 77512
rect 2459 77472 2504 77500
rect 2498 77460 2504 77472
rect 2556 77460 2562 77512
rect 3970 77500 3976 77512
rect 3931 77472 3976 77500
rect 3970 77460 3976 77472
rect 4028 77460 4034 77512
rect 4062 77460 4068 77512
rect 4120 77500 4126 77512
rect 5276 77509 5304 77540
rect 4617 77503 4675 77509
rect 4617 77500 4629 77503
rect 4120 77472 4629 77500
rect 4120 77460 4126 77472
rect 4617 77469 4629 77472
rect 4663 77469 4675 77503
rect 4617 77463 4675 77469
rect 5261 77503 5319 77509
rect 5261 77469 5273 77503
rect 5307 77469 5319 77503
rect 9398 77500 9404 77512
rect 9359 77472 9404 77500
rect 5261 77463 5319 77469
rect 9398 77460 9404 77472
rect 9456 77460 9462 77512
rect 10134 77500 10140 77512
rect 10095 77472 10140 77500
rect 10134 77460 10140 77472
rect 10192 77460 10198 77512
rect 1118 77392 1124 77444
rect 1176 77432 1182 77444
rect 1765 77435 1823 77441
rect 1765 77432 1777 77435
rect 1176 77404 1777 77432
rect 1176 77392 1182 77404
rect 1765 77401 1777 77404
rect 1811 77401 1823 77435
rect 1765 77395 1823 77401
rect 1949 77435 2007 77441
rect 1949 77401 1961 77435
rect 1995 77432 2007 77435
rect 2958 77432 2964 77444
rect 1995 77404 2964 77432
rect 1995 77401 2007 77404
rect 1949 77395 2007 77401
rect 2958 77392 2964 77404
rect 3016 77392 3022 77444
rect 3050 77324 3056 77376
rect 3108 77364 3114 77376
rect 3789 77367 3847 77373
rect 3789 77364 3801 77367
rect 3108 77336 3801 77364
rect 3108 77324 3114 77336
rect 3789 77333 3801 77336
rect 3835 77333 3847 77367
rect 3789 77327 3847 77333
rect 4433 77367 4491 77373
rect 4433 77333 4445 77367
rect 4479 77364 4491 77367
rect 4614 77364 4620 77376
rect 4479 77336 4620 77364
rect 4479 77333 4491 77336
rect 4433 77327 4491 77333
rect 4614 77324 4620 77336
rect 4672 77324 4678 77376
rect 5074 77364 5080 77376
rect 5035 77336 5080 77364
rect 5074 77324 5080 77336
rect 5132 77324 5138 77376
rect 9953 77367 10011 77373
rect 9953 77333 9965 77367
rect 9999 77364 10011 77367
rect 11057 77367 11115 77373
rect 11057 77364 11069 77367
rect 9999 77336 11069 77364
rect 9999 77333 10011 77336
rect 9953 77327 10011 77333
rect 11057 77333 11069 77336
rect 11103 77333 11115 77367
rect 11057 77327 11115 77333
rect 1104 77274 10856 77296
rect 1104 77222 4213 77274
rect 4265 77222 4277 77274
rect 4329 77222 4341 77274
rect 4393 77222 4405 77274
rect 4457 77222 4469 77274
rect 4521 77222 7477 77274
rect 7529 77222 7541 77274
rect 7593 77222 7605 77274
rect 7657 77222 7669 77274
rect 7721 77222 7733 77274
rect 7785 77222 10856 77274
rect 1104 77200 10856 77222
rect 1394 77024 1400 77036
rect 1355 76996 1400 77024
rect 1394 76984 1400 76996
rect 1452 76984 1458 77036
rect 2038 77024 2044 77036
rect 1999 76996 2044 77024
rect 2038 76984 2044 76996
rect 2096 76984 2102 77036
rect 2685 77027 2743 77033
rect 2685 76993 2697 77027
rect 2731 77024 2743 77027
rect 2774 77024 2780 77036
rect 2731 76996 2780 77024
rect 2731 76993 2743 76996
rect 2685 76987 2743 76993
rect 2774 76984 2780 76996
rect 2832 76984 2838 77036
rect 3326 77024 3332 77036
rect 3287 76996 3332 77024
rect 3326 76984 3332 76996
rect 3384 76984 3390 77036
rect 4154 77024 4160 77036
rect 4115 76996 4160 77024
rect 4154 76984 4160 76996
rect 4212 76984 4218 77036
rect 10134 77024 10140 77036
rect 10095 76996 10140 77024
rect 10134 76984 10140 76996
rect 10192 76984 10198 77036
rect 2869 76891 2927 76897
rect 2869 76857 2881 76891
rect 2915 76888 2927 76891
rect 3418 76888 3424 76900
rect 2915 76860 3424 76888
rect 2915 76857 2927 76860
rect 2869 76851 2927 76857
rect 3418 76848 3424 76860
rect 3476 76848 3482 76900
rect 1578 76820 1584 76832
rect 1539 76792 1584 76820
rect 1578 76780 1584 76792
rect 1636 76780 1642 76832
rect 2222 76820 2228 76832
rect 2183 76792 2228 76820
rect 2222 76780 2228 76792
rect 2280 76780 2286 76832
rect 3510 76820 3516 76832
rect 3471 76792 3516 76820
rect 3510 76780 3516 76792
rect 3568 76780 3574 76832
rect 3970 76820 3976 76832
rect 3931 76792 3976 76820
rect 3970 76780 3976 76792
rect 4028 76780 4034 76832
rect 9858 76780 9864 76832
rect 9916 76820 9922 76832
rect 9953 76823 10011 76829
rect 9953 76820 9965 76823
rect 9916 76792 9965 76820
rect 9916 76780 9922 76792
rect 9953 76789 9965 76792
rect 9999 76789 10011 76823
rect 9953 76783 10011 76789
rect 1104 76730 10856 76752
rect 1104 76678 2582 76730
rect 2634 76678 2646 76730
rect 2698 76678 2710 76730
rect 2762 76678 2774 76730
rect 2826 76678 2838 76730
rect 2890 76678 5845 76730
rect 5897 76678 5909 76730
rect 5961 76678 5973 76730
rect 6025 76678 6037 76730
rect 6089 76678 6101 76730
rect 6153 76678 9109 76730
rect 9161 76678 9173 76730
rect 9225 76678 9237 76730
rect 9289 76678 9301 76730
rect 9353 76678 9365 76730
rect 9417 76678 10856 76730
rect 1104 76656 10856 76678
rect 1854 76576 1860 76628
rect 1912 76616 1918 76628
rect 5074 76616 5080 76628
rect 1912 76588 5080 76616
rect 1912 76576 1918 76588
rect 5074 76576 5080 76588
rect 5132 76576 5138 76628
rect 1210 76508 1216 76560
rect 1268 76548 1274 76560
rect 2225 76551 2283 76557
rect 2225 76548 2237 76551
rect 1268 76520 2237 76548
rect 1268 76508 1274 76520
rect 2225 76517 2237 76520
rect 2271 76517 2283 76551
rect 2225 76511 2283 76517
rect 2774 76508 2780 76560
rect 2832 76548 2838 76560
rect 3878 76548 3884 76560
rect 2832 76520 3884 76548
rect 2832 76508 2838 76520
rect 3878 76508 3884 76520
rect 3936 76508 3942 76560
rect 3970 76480 3976 76492
rect 1872 76452 3976 76480
rect 1670 76412 1676 76424
rect 1631 76384 1676 76412
rect 1670 76372 1676 76384
rect 1728 76372 1734 76424
rect 1872 76421 1900 76452
rect 3970 76440 3976 76452
rect 4028 76440 4034 76492
rect 2130 76421 2136 76424
rect 1857 76415 1915 76421
rect 1857 76381 1869 76415
rect 1903 76381 1915 76415
rect 2093 76415 2136 76421
rect 2093 76412 2105 76415
rect 2043 76384 2105 76412
rect 1857 76375 1915 76381
rect 2093 76381 2105 76384
rect 2188 76412 2194 76424
rect 2774 76412 2780 76424
rect 2188 76384 2780 76412
rect 2093 76375 2136 76381
rect 2130 76372 2136 76375
rect 2188 76372 2194 76384
rect 2774 76372 2780 76384
rect 2832 76372 2838 76424
rect 2958 76412 2964 76424
rect 2919 76384 2964 76412
rect 2958 76372 2964 76384
rect 3016 76372 3022 76424
rect 10137 76415 10195 76421
rect 10137 76381 10149 76415
rect 10183 76412 10195 76415
rect 10965 76415 11023 76421
rect 10965 76412 10977 76415
rect 10183 76384 10977 76412
rect 10183 76381 10195 76384
rect 10137 76375 10195 76381
rect 10965 76381 10977 76384
rect 11011 76381 11023 76415
rect 10965 76375 11023 76381
rect 1949 76347 2007 76353
rect 1949 76313 1961 76347
rect 1995 76344 2007 76347
rect 1995 76316 6914 76344
rect 1995 76313 2007 76316
rect 1949 76307 2007 76313
rect 2777 76279 2835 76285
rect 2777 76245 2789 76279
rect 2823 76276 2835 76279
rect 3142 76276 3148 76288
rect 2823 76248 3148 76276
rect 2823 76245 2835 76248
rect 2777 76239 2835 76245
rect 3142 76236 3148 76248
rect 3200 76236 3206 76288
rect 6886 76276 6914 76316
rect 9953 76279 10011 76285
rect 9953 76276 9965 76279
rect 6886 76248 9965 76276
rect 9953 76245 9965 76248
rect 9999 76245 10011 76279
rect 9953 76239 10011 76245
rect 1104 76186 10856 76208
rect 1104 76134 4213 76186
rect 4265 76134 4277 76186
rect 4329 76134 4341 76186
rect 4393 76134 4405 76186
rect 4457 76134 4469 76186
rect 4521 76134 7477 76186
rect 7529 76134 7541 76186
rect 7593 76134 7605 76186
rect 7657 76134 7669 76186
rect 7721 76134 7733 76186
rect 7785 76134 10856 76186
rect 1104 76112 10856 76134
rect 4706 76072 4712 76084
rect 2884 76044 4712 76072
rect 1854 76004 1860 76016
rect 1815 75976 1860 76004
rect 1854 75964 1860 75976
rect 1912 75964 1918 76016
rect 1949 76007 2007 76013
rect 1949 75973 1961 76007
rect 1995 76004 2007 76007
rect 1995 75976 2774 76004
rect 1995 75973 2007 75976
rect 1949 75967 2007 75973
rect 937 75939 995 75945
rect 937 75905 949 75939
rect 983 75936 995 75939
rect 1670 75936 1676 75948
rect 983 75908 1676 75936
rect 983 75905 995 75908
rect 937 75899 995 75905
rect 1670 75896 1676 75908
rect 1728 75896 1734 75948
rect 2130 75945 2136 75948
rect 2093 75939 2136 75945
rect 2093 75905 2105 75939
rect 2093 75899 2136 75905
rect 2130 75896 2136 75899
rect 2188 75896 2194 75948
rect 2746 75936 2774 75976
rect 2884 75936 2912 76044
rect 4706 76032 4712 76044
rect 4764 76032 4770 76084
rect 2746 75908 2912 75936
rect 2961 75939 3019 75945
rect 2961 75905 2973 75939
rect 3007 75936 3019 75939
rect 3602 75936 3608 75948
rect 3007 75908 3608 75936
rect 3007 75905 3019 75908
rect 2961 75899 3019 75905
rect 3602 75896 3608 75908
rect 3660 75896 3666 75948
rect 6362 75936 6368 75948
rect 3712 75908 6368 75936
rect 2225 75803 2283 75809
rect 2225 75769 2237 75803
rect 2271 75800 2283 75803
rect 3712 75800 3740 75908
rect 6362 75896 6368 75908
rect 6420 75896 6426 75948
rect 10137 75939 10195 75945
rect 10137 75905 10149 75939
rect 10183 75936 10195 75939
rect 10183 75908 10272 75936
rect 10183 75905 10195 75908
rect 10137 75899 10195 75905
rect 10244 75880 10272 75908
rect 10226 75828 10232 75880
rect 10284 75828 10290 75880
rect 2271 75772 3740 75800
rect 2271 75769 2283 75772
rect 2225 75763 2283 75769
rect 1762 75692 1768 75744
rect 1820 75732 1826 75744
rect 2777 75735 2835 75741
rect 2777 75732 2789 75735
rect 1820 75704 2789 75732
rect 1820 75692 1826 75704
rect 2777 75701 2789 75704
rect 2823 75701 2835 75735
rect 9950 75732 9956 75744
rect 9911 75704 9956 75732
rect 2777 75695 2835 75701
rect 9950 75692 9956 75704
rect 10008 75692 10014 75744
rect 1104 75642 10856 75664
rect 1104 75590 2582 75642
rect 2634 75590 2646 75642
rect 2698 75590 2710 75642
rect 2762 75590 2774 75642
rect 2826 75590 2838 75642
rect 2890 75590 5845 75642
rect 5897 75590 5909 75642
rect 5961 75590 5973 75642
rect 6025 75590 6037 75642
rect 6089 75590 6101 75642
rect 6153 75590 9109 75642
rect 9161 75590 9173 75642
rect 9225 75590 9237 75642
rect 9289 75590 9301 75642
rect 9353 75590 9365 75642
rect 9417 75590 10856 75642
rect 1104 75568 10856 75590
rect 382 75420 388 75472
rect 440 75460 446 75472
rect 2409 75463 2467 75469
rect 2409 75460 2421 75463
rect 440 75432 2421 75460
rect 440 75420 446 75432
rect 2409 75429 2421 75432
rect 2455 75429 2467 75463
rect 2409 75423 2467 75429
rect 1302 75284 1308 75336
rect 1360 75324 1366 75336
rect 2590 75333 2596 75336
rect 1397 75327 1455 75333
rect 1397 75324 1409 75327
rect 1360 75296 1409 75324
rect 1360 75284 1366 75296
rect 1397 75293 1409 75296
rect 1443 75293 1455 75327
rect 2588 75324 2596 75333
rect 2551 75296 2596 75324
rect 1397 75287 1455 75293
rect 2588 75287 2596 75296
rect 2590 75284 2596 75287
rect 2648 75284 2654 75336
rect 2685 75327 2743 75333
rect 2685 75293 2697 75327
rect 2731 75324 2743 75327
rect 2731 75296 2912 75324
rect 2731 75293 2743 75296
rect 2685 75287 2743 75293
rect 2777 75259 2835 75265
rect 2777 75225 2789 75259
rect 2823 75225 2835 75259
rect 2884 75256 2912 75296
rect 2958 75284 2964 75336
rect 3016 75324 3022 75336
rect 3970 75324 3976 75336
rect 3016 75296 3061 75324
rect 3931 75296 3976 75324
rect 3016 75284 3022 75296
rect 3970 75284 3976 75296
rect 4028 75284 4034 75336
rect 10134 75324 10140 75336
rect 10095 75296 10140 75324
rect 10134 75284 10140 75296
rect 10192 75284 10198 75336
rect 2884 75228 6914 75256
rect 2777 75219 2835 75225
rect 1581 75191 1639 75197
rect 1581 75157 1593 75191
rect 1627 75188 1639 75191
rect 1854 75188 1860 75200
rect 1627 75160 1860 75188
rect 1627 75157 1639 75160
rect 1581 75151 1639 75157
rect 1854 75148 1860 75160
rect 1912 75148 1918 75200
rect 2792 75188 2820 75219
rect 3050 75188 3056 75200
rect 2792 75160 3056 75188
rect 3050 75148 3056 75160
rect 3108 75148 3114 75200
rect 3786 75188 3792 75200
rect 3747 75160 3792 75188
rect 3786 75148 3792 75160
rect 3844 75148 3850 75200
rect 6886 75188 6914 75228
rect 9953 75191 10011 75197
rect 9953 75188 9965 75191
rect 6886 75160 9965 75188
rect 9953 75157 9965 75160
rect 9999 75157 10011 75191
rect 9953 75151 10011 75157
rect 1104 75098 10856 75120
rect 1104 75046 4213 75098
rect 4265 75046 4277 75098
rect 4329 75046 4341 75098
rect 4393 75046 4405 75098
rect 4457 75046 4469 75098
rect 4521 75046 7477 75098
rect 7529 75046 7541 75098
rect 7593 75046 7605 75098
rect 7657 75046 7669 75098
rect 7721 75046 7733 75098
rect 7785 75046 10856 75098
rect 1104 75024 10856 75046
rect 2866 74944 2872 74996
rect 2924 74984 2930 74996
rect 4614 74984 4620 74996
rect 2924 74956 4620 74984
rect 2924 74944 2930 74956
rect 4614 74944 4620 74956
rect 4672 74944 4678 74996
rect 937 74919 995 74925
rect 937 74885 949 74919
rect 983 74916 995 74919
rect 983 74888 3464 74916
rect 983 74885 995 74888
rect 937 74879 995 74885
rect 1394 74848 1400 74860
rect 1355 74820 1400 74848
rect 1394 74808 1400 74820
rect 1452 74808 1458 74860
rect 2590 74857 2596 74860
rect 2588 74848 2596 74857
rect 2551 74820 2596 74848
rect 2588 74811 2596 74820
rect 2590 74808 2596 74811
rect 2648 74808 2654 74860
rect 2685 74851 2743 74857
rect 2685 74817 2697 74851
rect 2731 74817 2743 74851
rect 2685 74811 2743 74817
rect 2777 74851 2835 74857
rect 2777 74817 2789 74851
rect 2823 74848 2835 74851
rect 2866 74848 2872 74860
rect 2823 74820 2872 74848
rect 2823 74817 2835 74820
rect 2777 74811 2835 74817
rect 2700 74780 2728 74811
rect 2866 74808 2872 74820
rect 2924 74808 2930 74860
rect 2958 74808 2964 74860
rect 3016 74848 3022 74860
rect 3326 74848 3332 74860
rect 3016 74820 3332 74848
rect 3016 74808 3022 74820
rect 3326 74808 3332 74820
rect 3384 74808 3390 74860
rect 3436 74857 3464 74888
rect 3510 74876 3516 74928
rect 3568 74916 3574 74928
rect 3605 74919 3663 74925
rect 3605 74916 3617 74919
rect 3568 74888 3617 74916
rect 3568 74876 3574 74888
rect 3605 74885 3617 74888
rect 3651 74885 3663 74919
rect 3605 74879 3663 74885
rect 3697 74919 3755 74925
rect 3697 74885 3709 74919
rect 3743 74916 3755 74919
rect 9858 74916 9864 74928
rect 3743 74888 9864 74916
rect 3743 74885 3755 74888
rect 3697 74879 3755 74885
rect 9858 74876 9864 74888
rect 9916 74876 9922 74928
rect 3878 74857 3884 74860
rect 3421 74851 3479 74857
rect 3421 74817 3433 74851
rect 3467 74817 3479 74851
rect 3421 74811 3479 74817
rect 3841 74851 3884 74857
rect 3841 74817 3853 74851
rect 3841 74811 3884 74817
rect 3878 74808 3884 74811
rect 3936 74808 3942 74860
rect 9950 74780 9956 74792
rect 2700 74752 9956 74780
rect 9950 74740 9956 74752
rect 10008 74740 10014 74792
rect 4614 74712 4620 74724
rect 3896 74684 4620 74712
rect 1581 74647 1639 74653
rect 1581 74613 1593 74647
rect 1627 74644 1639 74647
rect 1946 74644 1952 74656
rect 1627 74616 1952 74644
rect 1627 74613 1639 74616
rect 1581 74607 1639 74613
rect 1946 74604 1952 74616
rect 2004 74604 2010 74656
rect 2409 74647 2467 74653
rect 2409 74613 2421 74647
rect 2455 74644 2467 74647
rect 3896 74644 3924 74684
rect 4614 74672 4620 74684
rect 4672 74672 4678 74724
rect 2455 74616 3924 74644
rect 3973 74647 4031 74653
rect 2455 74613 2467 74616
rect 2409 74607 2467 74613
rect 3973 74613 3985 74647
rect 4019 74644 4031 74647
rect 8294 74644 8300 74656
rect 4019 74616 8300 74644
rect 4019 74613 4031 74616
rect 3973 74607 4031 74613
rect 8294 74604 8300 74616
rect 8352 74604 8358 74656
rect 1104 74554 10856 74576
rect 1104 74502 2582 74554
rect 2634 74502 2646 74554
rect 2698 74502 2710 74554
rect 2762 74502 2774 74554
rect 2826 74502 2838 74554
rect 2890 74502 5845 74554
rect 5897 74502 5909 74554
rect 5961 74502 5973 74554
rect 6025 74502 6037 74554
rect 6089 74502 6101 74554
rect 6153 74502 9109 74554
rect 9161 74502 9173 74554
rect 9225 74502 9237 74554
rect 9289 74502 9301 74554
rect 9353 74502 9365 74554
rect 9417 74502 10856 74554
rect 1104 74480 10856 74502
rect 3605 74443 3663 74449
rect 3605 74440 3617 74443
rect 1688 74412 3617 74440
rect 1397 74239 1455 74245
rect 1397 74205 1409 74239
rect 1443 74205 1455 74239
rect 1578 74236 1584 74248
rect 1539 74208 1584 74236
rect 1397 74199 1455 74205
rect 1412 74100 1440 74199
rect 1578 74196 1584 74208
rect 1636 74196 1642 74248
rect 1688 74245 1716 74412
rect 3605 74409 3617 74412
rect 3651 74409 3663 74443
rect 3605 74403 3663 74409
rect 1949 74375 2007 74381
rect 1949 74341 1961 74375
rect 1995 74341 2007 74375
rect 1949 74335 2007 74341
rect 2593 74375 2651 74381
rect 2593 74341 2605 74375
rect 2639 74372 2651 74375
rect 4890 74372 4896 74384
rect 2639 74344 4896 74372
rect 2639 74341 2651 74344
rect 2593 74335 2651 74341
rect 1964 74304 1992 74335
rect 4890 74332 4896 74344
rect 4948 74332 4954 74384
rect 11333 74307 11391 74313
rect 11333 74304 11345 74307
rect 1964 74276 11345 74304
rect 11333 74273 11345 74276
rect 11379 74273 11391 74307
rect 11333 74267 11391 74273
rect 1673 74239 1731 74245
rect 1673 74205 1685 74239
rect 1719 74205 1731 74239
rect 1673 74199 1731 74205
rect 1770 74239 1828 74245
rect 1770 74205 1782 74239
rect 1816 74205 1828 74239
rect 1770 74199 1828 74205
rect 1486 74128 1492 74180
rect 1544 74168 1550 74180
rect 1785 74168 1813 74199
rect 2498 74196 2504 74248
rect 2556 74236 2562 74248
rect 2774 74245 2780 74248
rect 2731 74239 2780 74245
rect 2731 74236 2743 74239
rect 2556 74208 2743 74236
rect 2556 74196 2562 74208
rect 2731 74205 2743 74208
rect 2777 74205 2780 74239
rect 2731 74199 2780 74205
rect 2774 74196 2780 74199
rect 2832 74196 2838 74248
rect 2869 74239 2927 74245
rect 2869 74205 2881 74239
rect 2915 74236 2927 74239
rect 3145 74239 3203 74245
rect 2915 74208 3096 74236
rect 2915 74205 2927 74208
rect 2869 74199 2927 74205
rect 1544 74140 1813 74168
rect 2961 74171 3019 74177
rect 1544 74128 1550 74140
rect 2961 74137 2973 74171
rect 3007 74137 3019 74171
rect 3068 74168 3096 74208
rect 3145 74205 3157 74239
rect 3191 74236 3203 74239
rect 3326 74236 3332 74248
rect 3191 74208 3332 74236
rect 3191 74205 3203 74208
rect 3145 74199 3203 74205
rect 3326 74196 3332 74208
rect 3384 74196 3390 74248
rect 10134 74236 10140 74248
rect 10095 74208 10140 74236
rect 10134 74196 10140 74208
rect 10192 74196 10198 74248
rect 3068 74140 9996 74168
rect 2961 74131 3019 74137
rect 2130 74100 2136 74112
rect 1412 74072 2136 74100
rect 2130 74060 2136 74072
rect 2188 74060 2194 74112
rect 2976 74100 3004 74131
rect 3234 74100 3240 74112
rect 2976 74072 3240 74100
rect 3234 74060 3240 74072
rect 3292 74060 3298 74112
rect 3605 74103 3663 74109
rect 3605 74069 3617 74103
rect 3651 74100 3663 74103
rect 9766 74100 9772 74112
rect 3651 74072 9772 74100
rect 3651 74069 3663 74072
rect 3605 74063 3663 74069
rect 9766 74060 9772 74072
rect 9824 74060 9830 74112
rect 9968 74109 9996 74140
rect 9953 74103 10011 74109
rect 9953 74069 9965 74103
rect 9999 74069 10011 74103
rect 9953 74063 10011 74069
rect 1104 74010 10856 74032
rect 1104 73958 4213 74010
rect 4265 73958 4277 74010
rect 4329 73958 4341 74010
rect 4393 73958 4405 74010
rect 4457 73958 4469 74010
rect 4521 73958 7477 74010
rect 7529 73958 7541 74010
rect 7593 73958 7605 74010
rect 7657 73958 7669 74010
rect 7721 73958 7733 74010
rect 7785 73958 10856 74010
rect 1104 73936 10856 73958
rect 1857 73831 1915 73837
rect 1857 73797 1869 73831
rect 1903 73828 1915 73831
rect 3142 73828 3148 73840
rect 1903 73800 3148 73828
rect 1903 73797 1915 73800
rect 1857 73791 1915 73797
rect 3142 73788 3148 73800
rect 3200 73788 3206 73840
rect 1486 73720 1492 73772
rect 1544 73760 1550 73772
rect 1621 73763 1679 73769
rect 1621 73760 1633 73763
rect 1544 73732 1633 73760
rect 1544 73720 1550 73732
rect 1621 73729 1633 73732
rect 1667 73729 1679 73763
rect 1621 73723 1679 73729
rect 1765 73763 1823 73769
rect 1765 73729 1777 73763
rect 1811 73729 1823 73763
rect 1765 73723 1823 73729
rect 2041 73763 2099 73769
rect 2041 73729 2053 73763
rect 2087 73760 2099 73763
rect 2130 73760 2136 73772
rect 2087 73732 2136 73760
rect 2087 73729 2099 73732
rect 2041 73723 2099 73729
rect 1780 73692 1808 73723
rect 2130 73720 2136 73732
rect 2188 73720 2194 73772
rect 2685 73763 2743 73769
rect 2685 73729 2697 73763
rect 2731 73760 2743 73763
rect 2958 73760 2964 73772
rect 2731 73732 2964 73760
rect 2731 73729 2743 73732
rect 2685 73723 2743 73729
rect 2958 73720 2964 73732
rect 3016 73720 3022 73772
rect 10134 73760 10140 73772
rect 10095 73732 10140 73760
rect 10134 73720 10140 73732
rect 10192 73720 10198 73772
rect 9950 73692 9956 73704
rect 1780 73664 9956 73692
rect 9950 73652 9956 73664
rect 10008 73652 10014 73704
rect 1489 73627 1547 73633
rect 1489 73593 1501 73627
rect 1535 73624 1547 73627
rect 5534 73624 5540 73636
rect 1535 73596 5540 73624
rect 1535 73593 1547 73596
rect 1489 73587 1547 73593
rect 5534 73584 5540 73596
rect 5592 73584 5598 73636
rect 2314 73516 2320 73568
rect 2372 73556 2378 73568
rect 2501 73559 2559 73565
rect 2501 73556 2513 73559
rect 2372 73528 2513 73556
rect 2372 73516 2378 73528
rect 2501 73525 2513 73528
rect 2547 73525 2559 73559
rect 2501 73519 2559 73525
rect 9953 73559 10011 73565
rect 9953 73525 9965 73559
rect 9999 73556 10011 73559
rect 11057 73559 11115 73565
rect 11057 73556 11069 73559
rect 9999 73528 11069 73556
rect 9999 73525 10011 73528
rect 9953 73519 10011 73525
rect 11057 73525 11069 73528
rect 11103 73525 11115 73559
rect 11057 73519 11115 73525
rect 1104 73466 10856 73488
rect 1104 73414 2582 73466
rect 2634 73414 2646 73466
rect 2698 73414 2710 73466
rect 2762 73414 2774 73466
rect 2826 73414 2838 73466
rect 2890 73414 5845 73466
rect 5897 73414 5909 73466
rect 5961 73414 5973 73466
rect 6025 73414 6037 73466
rect 6089 73414 6101 73466
rect 6153 73414 9109 73466
rect 9161 73414 9173 73466
rect 9225 73414 9237 73466
rect 9289 73414 9301 73466
rect 9353 73414 9365 73466
rect 9417 73414 10856 73466
rect 1104 73392 10856 73414
rect 1394 73148 1400 73160
rect 1355 73120 1400 73148
rect 1394 73108 1400 73120
rect 1452 73108 1458 73160
rect 2222 73148 2228 73160
rect 2183 73120 2228 73148
rect 2222 73108 2228 73120
rect 2280 73108 2286 73160
rect 10134 73148 10140 73160
rect 10095 73120 10140 73148
rect 10134 73108 10140 73120
rect 10192 73108 10198 73160
rect 1581 73015 1639 73021
rect 1581 72981 1593 73015
rect 1627 73012 1639 73015
rect 1670 73012 1676 73024
rect 1627 72984 1676 73012
rect 1627 72981 1639 72984
rect 1581 72975 1639 72981
rect 1670 72972 1676 72984
rect 1728 72972 1734 73024
rect 2038 73012 2044 73024
rect 1999 72984 2044 73012
rect 2038 72972 2044 72984
rect 2096 72972 2102 73024
rect 9953 73015 10011 73021
rect 9953 72981 9965 73015
rect 9999 73012 10011 73015
rect 11149 73015 11207 73021
rect 11149 73012 11161 73015
rect 9999 72984 11161 73012
rect 9999 72981 10011 72984
rect 9953 72975 10011 72981
rect 11149 72981 11161 72984
rect 11195 72981 11207 73015
rect 11149 72975 11207 72981
rect 1104 72922 10856 72944
rect 1104 72870 4213 72922
rect 4265 72870 4277 72922
rect 4329 72870 4341 72922
rect 4393 72870 4405 72922
rect 4457 72870 4469 72922
rect 4521 72870 7477 72922
rect 7529 72870 7541 72922
rect 7593 72870 7605 72922
rect 7657 72870 7669 72922
rect 7721 72870 7733 72922
rect 7785 72870 10856 72922
rect 1104 72848 10856 72870
rect 1302 72632 1308 72684
rect 1360 72672 1366 72684
rect 1397 72675 1455 72681
rect 1397 72672 1409 72675
rect 1360 72644 1409 72672
rect 1360 72632 1366 72644
rect 1397 72641 1409 72644
rect 1443 72641 1455 72675
rect 1397 72635 1455 72641
rect 1581 72471 1639 72477
rect 1581 72437 1593 72471
rect 1627 72468 1639 72471
rect 2222 72468 2228 72480
rect 1627 72440 2228 72468
rect 1627 72437 1639 72440
rect 1581 72431 1639 72437
rect 2222 72428 2228 72440
rect 2280 72428 2286 72480
rect 1104 72378 10856 72400
rect 1104 72326 2582 72378
rect 2634 72326 2646 72378
rect 2698 72326 2710 72378
rect 2762 72326 2774 72378
rect 2826 72326 2838 72378
rect 2890 72326 5845 72378
rect 5897 72326 5909 72378
rect 5961 72326 5973 72378
rect 6025 72326 6037 72378
rect 6089 72326 6101 72378
rect 6153 72326 9109 72378
rect 9161 72326 9173 72378
rect 9225 72326 9237 72378
rect 9289 72326 9301 72378
rect 9353 72326 9365 72378
rect 9417 72326 10856 72378
rect 1104 72304 10856 72326
rect 1394 72224 1400 72276
rect 1452 72264 1458 72276
rect 2130 72264 2136 72276
rect 1452 72236 2136 72264
rect 1452 72224 1458 72236
rect 2130 72224 2136 72236
rect 2188 72224 2194 72276
rect 9950 72264 9956 72276
rect 9911 72236 9956 72264
rect 9950 72224 9956 72236
rect 10008 72224 10014 72276
rect 1949 72199 2007 72205
rect 1949 72165 1961 72199
rect 1995 72196 2007 72199
rect 11241 72199 11299 72205
rect 11241 72196 11253 72199
rect 1995 72168 11253 72196
rect 1995 72165 2007 72168
rect 1949 72159 2007 72165
rect 11241 72165 11253 72168
rect 11287 72165 11299 72199
rect 11241 72159 11299 72165
rect 3786 72128 3792 72140
rect 1596 72100 3792 72128
rect 1394 72060 1400 72072
rect 1355 72032 1400 72060
rect 1394 72020 1400 72032
rect 1452 72020 1458 72072
rect 1596 72069 1624 72100
rect 3786 72088 3792 72100
rect 3844 72088 3850 72140
rect 1581 72063 1639 72069
rect 1581 72029 1593 72063
rect 1627 72029 1639 72063
rect 1762 72060 1768 72072
rect 1727 72032 1768 72060
rect 1581 72023 1639 72029
rect 1762 72020 1768 72032
rect 1820 72069 1826 72072
rect 1820 72063 1875 72069
rect 1820 72029 1829 72063
rect 1863 72060 1875 72063
rect 3234 72060 3240 72072
rect 1863 72032 3240 72060
rect 1863 72029 1875 72032
rect 1820 72023 1875 72029
rect 1820 72020 1826 72023
rect 3234 72020 3240 72032
rect 3292 72020 3298 72072
rect 10134 72060 10140 72072
rect 10095 72032 10140 72060
rect 10134 72020 10140 72032
rect 10192 72020 10198 72072
rect 1673 71995 1731 72001
rect 1673 71961 1685 71995
rect 1719 71992 1731 71995
rect 9858 71992 9864 72004
rect 1719 71964 9864 71992
rect 1719 71961 1731 71964
rect 1673 71955 1731 71961
rect 9858 71952 9864 71964
rect 9916 71952 9922 72004
rect 1486 71884 1492 71936
rect 1544 71924 1550 71936
rect 1762 71924 1768 71936
rect 1544 71896 1768 71924
rect 1544 71884 1550 71896
rect 1762 71884 1768 71896
rect 1820 71884 1826 71936
rect 1104 71834 10856 71856
rect 1104 71782 4213 71834
rect 4265 71782 4277 71834
rect 4329 71782 4341 71834
rect 4393 71782 4405 71834
rect 4457 71782 4469 71834
rect 4521 71782 7477 71834
rect 7529 71782 7541 71834
rect 7593 71782 7605 71834
rect 7657 71782 7669 71834
rect 7721 71782 7733 71834
rect 7785 71782 10856 71834
rect 1104 71760 10856 71782
rect 9766 71680 9772 71732
rect 9824 71720 9830 71732
rect 9953 71723 10011 71729
rect 9953 71720 9965 71723
rect 9824 71692 9965 71720
rect 9824 71680 9830 71692
rect 9953 71689 9965 71692
rect 9999 71689 10011 71723
rect 9953 71683 10011 71689
rect 10134 71584 10140 71596
rect 10095 71556 10140 71584
rect 10134 71544 10140 71556
rect 10192 71544 10198 71596
rect 1394 71516 1400 71528
rect 1355 71488 1400 71516
rect 1394 71476 1400 71488
rect 1452 71476 1458 71528
rect 1673 71519 1731 71525
rect 1673 71485 1685 71519
rect 1719 71516 1731 71519
rect 1762 71516 1768 71528
rect 1719 71488 1768 71516
rect 1719 71485 1731 71488
rect 1673 71479 1731 71485
rect 1762 71476 1768 71488
rect 1820 71476 1826 71528
rect 1104 71290 10856 71312
rect 1104 71238 2582 71290
rect 2634 71238 2646 71290
rect 2698 71238 2710 71290
rect 2762 71238 2774 71290
rect 2826 71238 2838 71290
rect 2890 71238 5845 71290
rect 5897 71238 5909 71290
rect 5961 71238 5973 71290
rect 6025 71238 6037 71290
rect 6089 71238 6101 71290
rect 6153 71238 9109 71290
rect 9161 71238 9173 71290
rect 9225 71238 9237 71290
rect 9289 71238 9301 71290
rect 9353 71238 9365 71290
rect 9417 71238 10856 71290
rect 1104 71216 10856 71238
rect 1302 71000 1308 71052
rect 1360 71040 1366 71052
rect 1397 71043 1455 71049
rect 1397 71040 1409 71043
rect 1360 71012 1409 71040
rect 1360 71000 1366 71012
rect 1397 71009 1409 71012
rect 1443 71009 1455 71043
rect 1397 71003 1455 71009
rect 1673 70975 1731 70981
rect 1673 70941 1685 70975
rect 1719 70972 1731 70975
rect 2498 70972 2504 70984
rect 1719 70944 2504 70972
rect 1719 70941 1731 70944
rect 1673 70935 1731 70941
rect 2498 70932 2504 70944
rect 2556 70932 2562 70984
rect 2685 70975 2743 70981
rect 2685 70941 2697 70975
rect 2731 70972 2743 70975
rect 2774 70972 2780 70984
rect 2731 70944 2780 70972
rect 2731 70941 2743 70944
rect 2685 70935 2743 70941
rect 2774 70932 2780 70944
rect 2832 70932 2838 70984
rect 2869 70839 2927 70845
rect 2869 70805 2881 70839
rect 2915 70836 2927 70839
rect 4062 70836 4068 70848
rect 2915 70808 4068 70836
rect 2915 70805 2927 70808
rect 2869 70799 2927 70805
rect 4062 70796 4068 70808
rect 4120 70796 4126 70848
rect 1104 70746 10856 70768
rect 1104 70694 4213 70746
rect 4265 70694 4277 70746
rect 4329 70694 4341 70746
rect 4393 70694 4405 70746
rect 4457 70694 4469 70746
rect 4521 70694 7477 70746
rect 7529 70694 7541 70746
rect 7593 70694 7605 70746
rect 7657 70694 7669 70746
rect 7721 70694 7733 70746
rect 7785 70694 10856 70746
rect 1104 70672 10856 70694
rect 2682 70632 2688 70644
rect 1688 70604 2688 70632
rect 1688 70573 1716 70604
rect 2682 70592 2688 70604
rect 2740 70592 2746 70644
rect 2866 70592 2872 70644
rect 2924 70632 2930 70644
rect 3418 70632 3424 70644
rect 2924 70604 3424 70632
rect 2924 70592 2930 70604
rect 3418 70592 3424 70604
rect 3476 70592 3482 70644
rect 9858 70592 9864 70644
rect 9916 70632 9922 70644
rect 9953 70635 10011 70641
rect 9953 70632 9965 70635
rect 9916 70604 9965 70632
rect 9916 70592 9922 70604
rect 9953 70601 9965 70604
rect 9999 70601 10011 70635
rect 9953 70595 10011 70601
rect 1673 70567 1731 70573
rect 1673 70533 1685 70567
rect 1719 70533 1731 70567
rect 1673 70527 1731 70533
rect 2593 70567 2651 70573
rect 2593 70533 2605 70567
rect 2639 70564 2651 70567
rect 11057 70567 11115 70573
rect 11057 70564 11069 70567
rect 2639 70536 11069 70564
rect 2639 70533 2651 70536
rect 2593 70527 2651 70533
rect 11057 70533 11069 70536
rect 11103 70533 11115 70567
rect 11057 70527 11115 70533
rect 2449 70499 2507 70505
rect 2449 70496 2461 70499
rect 2240 70468 2461 70496
rect 934 70320 940 70372
rect 992 70360 998 70372
rect 1762 70360 1768 70372
rect 992 70332 1768 70360
rect 992 70320 998 70332
rect 1762 70320 1768 70332
rect 1820 70320 1826 70372
rect 1578 70292 1584 70304
rect 1539 70264 1584 70292
rect 1578 70252 1584 70264
rect 1636 70252 1642 70304
rect 2240 70292 2268 70468
rect 2449 70465 2461 70468
rect 2495 70465 2507 70499
rect 2449 70459 2507 70465
rect 2685 70499 2743 70505
rect 2685 70465 2697 70499
rect 2731 70496 2743 70499
rect 2774 70496 2780 70508
rect 2731 70468 2780 70496
rect 2731 70465 2743 70468
rect 2685 70459 2743 70465
rect 2774 70456 2780 70468
rect 2832 70456 2838 70508
rect 2869 70499 2927 70505
rect 2869 70465 2881 70499
rect 2915 70496 2927 70499
rect 2958 70496 2964 70508
rect 2915 70468 2964 70496
rect 2915 70465 2927 70468
rect 2869 70459 2927 70465
rect 2958 70456 2964 70468
rect 3016 70496 3022 70508
rect 3326 70496 3332 70508
rect 3016 70468 3332 70496
rect 3016 70456 3022 70468
rect 3326 70456 3332 70468
rect 3384 70456 3390 70508
rect 3510 70496 3516 70508
rect 3471 70468 3516 70496
rect 3510 70456 3516 70468
rect 3568 70456 3574 70508
rect 10134 70496 10140 70508
rect 10095 70468 10140 70496
rect 10134 70456 10140 70468
rect 10192 70456 10198 70508
rect 7006 70428 7012 70440
rect 2332 70400 7012 70428
rect 2332 70369 2360 70400
rect 7006 70388 7012 70400
rect 7064 70388 7070 70440
rect 11057 70431 11115 70437
rect 11057 70397 11069 70431
rect 11103 70428 11115 70431
rect 11333 70431 11391 70437
rect 11333 70428 11345 70431
rect 11103 70400 11345 70428
rect 11103 70397 11115 70400
rect 11057 70391 11115 70397
rect 11333 70397 11345 70400
rect 11379 70397 11391 70431
rect 11333 70391 11391 70397
rect 2317 70363 2375 70369
rect 2317 70329 2329 70363
rect 2363 70360 2375 70363
rect 2363 70332 2397 70360
rect 2363 70329 2375 70332
rect 2317 70323 2375 70329
rect 2774 70320 2780 70372
rect 2832 70360 2838 70372
rect 3142 70360 3148 70372
rect 2832 70332 3148 70360
rect 2832 70320 2838 70332
rect 3142 70320 3148 70332
rect 3200 70320 3206 70372
rect 3050 70292 3056 70304
rect 2240 70264 3056 70292
rect 3050 70252 3056 70264
rect 3108 70252 3114 70304
rect 3329 70295 3387 70301
rect 3329 70261 3341 70295
rect 3375 70292 3387 70295
rect 3602 70292 3608 70304
rect 3375 70264 3608 70292
rect 3375 70261 3387 70264
rect 3329 70255 3387 70261
rect 3602 70252 3608 70264
rect 3660 70252 3666 70304
rect 1104 70202 10856 70224
rect 1104 70150 2582 70202
rect 2634 70150 2646 70202
rect 2698 70150 2710 70202
rect 2762 70150 2774 70202
rect 2826 70150 2838 70202
rect 2890 70150 5845 70202
rect 5897 70150 5909 70202
rect 5961 70150 5973 70202
rect 6025 70150 6037 70202
rect 6089 70150 6101 70202
rect 6153 70150 9109 70202
rect 9161 70150 9173 70202
rect 9225 70150 9237 70202
rect 9289 70150 9301 70202
rect 9353 70150 9365 70202
rect 9417 70150 10856 70202
rect 1104 70128 10856 70150
rect 2409 70023 2467 70029
rect 2409 69989 2421 70023
rect 2455 70020 2467 70023
rect 11793 70023 11851 70029
rect 11793 70020 11805 70023
rect 2455 69992 11805 70020
rect 2455 69989 2467 69992
rect 2409 69983 2467 69989
rect 11793 69989 11805 69992
rect 11839 69989 11851 70023
rect 11793 69983 11851 69989
rect 2866 69952 2872 69964
rect 2608 69924 2872 69952
rect 1302 69844 1308 69896
rect 1360 69884 1366 69896
rect 2608 69893 2636 69924
rect 2866 69912 2872 69924
rect 2924 69952 2930 69964
rect 3050 69952 3056 69964
rect 2924 69924 3056 69952
rect 2924 69912 2930 69924
rect 3050 69912 3056 69924
rect 3108 69912 3114 69964
rect 1397 69887 1455 69893
rect 1397 69884 1409 69887
rect 1360 69856 1409 69884
rect 1360 69844 1366 69856
rect 1397 69853 1409 69856
rect 1443 69853 1455 69887
rect 1397 69847 1455 69853
rect 2588 69887 2646 69893
rect 2588 69853 2600 69887
rect 2634 69853 2646 69887
rect 2588 69847 2646 69853
rect 2685 69887 2743 69893
rect 2685 69853 2697 69887
rect 2731 69884 2743 69887
rect 2961 69887 3019 69893
rect 2731 69856 2912 69884
rect 2731 69853 2743 69856
rect 2685 69847 2743 69853
rect 2406 69776 2412 69828
rect 2464 69816 2470 69828
rect 2777 69819 2835 69825
rect 2777 69816 2789 69819
rect 2464 69788 2789 69816
rect 2464 69776 2470 69788
rect 2777 69785 2789 69788
rect 2823 69785 2835 69819
rect 2884 69816 2912 69856
rect 2961 69853 2973 69887
rect 3007 69884 3019 69887
rect 3234 69884 3240 69896
rect 3007 69856 3240 69884
rect 3007 69853 3019 69856
rect 2961 69847 3019 69853
rect 3234 69844 3240 69856
rect 3292 69844 3298 69896
rect 3970 69884 3976 69896
rect 3931 69856 3976 69884
rect 3970 69844 3976 69856
rect 4028 69844 4034 69896
rect 10134 69884 10140 69896
rect 10095 69856 10140 69884
rect 10134 69844 10140 69856
rect 10192 69844 10198 69896
rect 11149 69819 11207 69825
rect 11149 69816 11161 69819
rect 2884 69788 11161 69816
rect 2777 69779 2835 69785
rect 11149 69785 11161 69788
rect 11195 69785 11207 69819
rect 11149 69779 11207 69785
rect 1581 69751 1639 69757
rect 1581 69717 1593 69751
rect 1627 69748 1639 69751
rect 3510 69748 3516 69760
rect 1627 69720 3516 69748
rect 1627 69717 1639 69720
rect 1581 69711 1639 69717
rect 3510 69708 3516 69720
rect 3568 69708 3574 69760
rect 3694 69708 3700 69760
rect 3752 69748 3758 69760
rect 3789 69751 3847 69757
rect 3789 69748 3801 69751
rect 3752 69720 3801 69748
rect 3752 69708 3758 69720
rect 3789 69717 3801 69720
rect 3835 69717 3847 69751
rect 9950 69748 9956 69760
rect 9911 69720 9956 69748
rect 3789 69711 3847 69717
rect 9950 69708 9956 69720
rect 10008 69708 10014 69760
rect 1104 69658 10856 69680
rect 1104 69606 4213 69658
rect 4265 69606 4277 69658
rect 4329 69606 4341 69658
rect 4393 69606 4405 69658
rect 4457 69606 4469 69658
rect 4521 69606 7477 69658
rect 7529 69606 7541 69658
rect 7593 69606 7605 69658
rect 7657 69606 7669 69658
rect 7721 69606 7733 69658
rect 7785 69606 10856 69658
rect 1104 69584 10856 69606
rect 1578 69504 1584 69556
rect 1636 69544 1642 69556
rect 3326 69544 3332 69556
rect 1636 69516 3332 69544
rect 1636 69504 1642 69516
rect 3326 69504 3332 69516
rect 3384 69504 3390 69556
rect 1762 69476 1768 69488
rect 1723 69448 1768 69476
rect 1762 69436 1768 69448
rect 1820 69436 1826 69488
rect 2130 69476 2136 69488
rect 1964 69448 2136 69476
rect 1578 69368 1584 69420
rect 1636 69417 1642 69420
rect 1636 69411 1685 69417
rect 1636 69377 1639 69411
rect 1673 69377 1685 69411
rect 1636 69371 1685 69377
rect 1857 69411 1915 69417
rect 1857 69377 1869 69411
rect 1903 69408 1915 69411
rect 1964 69408 1992 69448
rect 2130 69436 2136 69448
rect 2188 69436 2194 69488
rect 5718 69436 5724 69488
rect 5776 69476 5782 69488
rect 9950 69476 9956 69488
rect 5776 69448 9956 69476
rect 5776 69436 5782 69448
rect 9950 69436 9956 69448
rect 10008 69436 10014 69488
rect 1903 69380 1992 69408
rect 2041 69411 2099 69417
rect 1903 69377 1915 69380
rect 1857 69371 1915 69377
rect 2041 69377 2053 69411
rect 2087 69408 2099 69411
rect 2406 69408 2412 69420
rect 2087 69380 2412 69408
rect 2087 69377 2099 69380
rect 2041 69371 2099 69377
rect 1636 69368 1642 69371
rect 2406 69368 2412 69380
rect 2464 69368 2470 69420
rect 2958 69368 2964 69420
rect 3016 69408 3022 69420
rect 3053 69411 3111 69417
rect 3053 69408 3065 69411
rect 3016 69380 3065 69408
rect 3016 69368 3022 69380
rect 3053 69377 3065 69380
rect 3099 69408 3111 69411
rect 3234 69408 3240 69420
rect 3099 69380 3240 69408
rect 3099 69377 3111 69380
rect 3053 69371 3111 69377
rect 3234 69368 3240 69380
rect 3292 69368 3298 69420
rect 4154 69368 4160 69420
rect 4212 69408 4218 69420
rect 4249 69411 4307 69417
rect 4249 69408 4261 69411
rect 4212 69380 4261 69408
rect 4212 69368 4218 69380
rect 4249 69377 4261 69380
rect 4295 69377 4307 69411
rect 10134 69408 10140 69420
rect 10095 69380 10140 69408
rect 4249 69371 4307 69377
rect 10134 69368 10140 69380
rect 10192 69368 10198 69420
rect 937 69343 995 69349
rect 937 69309 949 69343
rect 983 69340 995 69343
rect 1762 69340 1768 69352
rect 983 69312 1768 69340
rect 983 69309 995 69312
rect 937 69303 995 69309
rect 1762 69300 1768 69312
rect 1820 69300 1826 69352
rect 2777 69343 2835 69349
rect 2777 69309 2789 69343
rect 2823 69340 2835 69343
rect 3142 69340 3148 69352
rect 2823 69312 3148 69340
rect 2823 69309 2835 69312
rect 2777 69303 2835 69309
rect 3142 69300 3148 69312
rect 3200 69300 3206 69352
rect 1394 69232 1400 69284
rect 1452 69272 1458 69284
rect 4065 69275 4123 69281
rect 4065 69272 4077 69275
rect 1452 69244 4077 69272
rect 1452 69232 1458 69244
rect 4065 69241 4077 69244
rect 4111 69241 4123 69275
rect 4065 69235 4123 69241
rect 1486 69204 1492 69216
rect 1447 69176 1492 69204
rect 1486 69164 1492 69176
rect 1544 69164 1550 69216
rect 9950 69204 9956 69216
rect 9911 69176 9956 69204
rect 9950 69164 9956 69176
rect 10008 69164 10014 69216
rect 1104 69114 10856 69136
rect 1104 69062 2582 69114
rect 2634 69062 2646 69114
rect 2698 69062 2710 69114
rect 2762 69062 2774 69114
rect 2826 69062 2838 69114
rect 2890 69062 5845 69114
rect 5897 69062 5909 69114
rect 5961 69062 5973 69114
rect 6025 69062 6037 69114
rect 6089 69062 6101 69114
rect 6153 69062 9109 69114
rect 9161 69062 9173 69114
rect 9225 69062 9237 69114
rect 9289 69062 9301 69114
rect 9353 69062 9365 69114
rect 9417 69062 10856 69114
rect 1104 69040 10856 69062
rect 2958 68864 2964 68876
rect 2919 68836 2964 68864
rect 2958 68824 2964 68836
rect 3016 68824 3022 68876
rect 1302 68756 1308 68808
rect 1360 68796 1366 68808
rect 1397 68799 1455 68805
rect 1397 68796 1409 68799
rect 1360 68768 1409 68796
rect 1360 68756 1366 68768
rect 1397 68765 1409 68768
rect 1443 68765 1455 68799
rect 1397 68759 1455 68765
rect 3237 68799 3295 68805
rect 3237 68765 3249 68799
rect 3283 68765 3295 68799
rect 3970 68796 3976 68808
rect 3931 68768 3976 68796
rect 3237 68759 3295 68765
rect 2958 68688 2964 68740
rect 3016 68728 3022 68740
rect 3252 68728 3280 68759
rect 3970 68756 3976 68768
rect 4028 68756 4034 68808
rect 3016 68700 3280 68728
rect 3016 68688 3022 68700
rect 1581 68663 1639 68669
rect 1581 68629 1593 68663
rect 1627 68660 1639 68663
rect 2130 68660 2136 68672
rect 1627 68632 2136 68660
rect 1627 68629 1639 68632
rect 1581 68623 1639 68629
rect 2130 68620 2136 68632
rect 2188 68620 2194 68672
rect 3786 68660 3792 68672
rect 3747 68632 3792 68660
rect 3786 68620 3792 68632
rect 3844 68620 3850 68672
rect 1104 68570 10856 68592
rect 1104 68518 4213 68570
rect 4265 68518 4277 68570
rect 4329 68518 4341 68570
rect 4393 68518 4405 68570
rect 4457 68518 4469 68570
rect 4521 68518 7477 68570
rect 7529 68518 7541 68570
rect 7593 68518 7605 68570
rect 7657 68518 7669 68570
rect 7721 68518 7733 68570
rect 7785 68518 10856 68570
rect 1104 68496 10856 68518
rect 1854 68416 1860 68468
rect 1912 68456 1918 68468
rect 1912 68428 3096 68456
rect 1912 68416 1918 68428
rect 1946 68388 1952 68400
rect 1907 68360 1952 68388
rect 1946 68348 1952 68360
rect 2004 68348 2010 68400
rect 3068 68397 3096 68428
rect 3234 68416 3240 68468
rect 3292 68456 3298 68468
rect 3973 68459 4031 68465
rect 3973 68456 3985 68459
rect 3292 68428 3985 68456
rect 3292 68416 3298 68428
rect 3973 68425 3985 68428
rect 4019 68425 4031 68459
rect 3973 68419 4031 68425
rect 2041 68391 2099 68397
rect 2041 68357 2053 68391
rect 2087 68388 2099 68391
rect 3053 68391 3111 68397
rect 2087 68360 2268 68388
rect 2087 68357 2099 68360
rect 2041 68351 2099 68357
rect 1670 68280 1676 68332
rect 1728 68320 1734 68332
rect 1765 68323 1823 68329
rect 1765 68320 1777 68323
rect 1728 68292 1777 68320
rect 1728 68280 1734 68292
rect 1765 68289 1777 68292
rect 1811 68289 1823 68323
rect 1765 68283 1823 68289
rect 2138 68323 2196 68329
rect 2138 68289 2150 68323
rect 2184 68289 2196 68323
rect 2138 68283 2196 68289
rect 1486 68212 1492 68264
rect 1544 68252 1550 68264
rect 2148 68252 2176 68283
rect 1544 68224 2176 68252
rect 1544 68212 1550 68224
rect 2240 68116 2268 68360
rect 3053 68357 3065 68391
rect 3099 68357 3111 68391
rect 3053 68351 3111 68357
rect 3145 68391 3203 68397
rect 3145 68357 3157 68391
rect 3191 68388 3203 68391
rect 9950 68388 9956 68400
rect 3191 68360 9956 68388
rect 3191 68357 3203 68360
rect 3145 68351 3203 68357
rect 9950 68348 9956 68360
rect 10008 68348 10014 68400
rect 2406 68280 2412 68332
rect 2464 68320 2470 68332
rect 3326 68329 3332 68332
rect 2869 68323 2927 68329
rect 2869 68320 2881 68323
rect 2464 68292 2881 68320
rect 2464 68280 2470 68292
rect 2869 68289 2881 68292
rect 2915 68289 2927 68323
rect 2869 68283 2927 68289
rect 3289 68323 3332 68329
rect 3289 68289 3301 68323
rect 3289 68283 3332 68289
rect 3326 68280 3332 68283
rect 3384 68280 3390 68332
rect 3418 68280 3424 68332
rect 3476 68320 3482 68332
rect 4157 68323 4215 68329
rect 4157 68320 4169 68323
rect 3476 68292 4169 68320
rect 3476 68280 3482 68292
rect 4157 68289 4169 68292
rect 4203 68289 4215 68323
rect 10134 68320 10140 68332
rect 10095 68292 10140 68320
rect 4157 68283 4215 68289
rect 10134 68280 10140 68292
rect 10192 68280 10198 68332
rect 7098 68252 7104 68264
rect 2746 68224 7104 68252
rect 2317 68187 2375 68193
rect 2317 68153 2329 68187
rect 2363 68184 2375 68187
rect 2746 68184 2774 68224
rect 7098 68212 7104 68224
rect 7156 68212 7162 68264
rect 9953 68187 10011 68193
rect 9953 68184 9965 68187
rect 2363 68156 2774 68184
rect 3344 68156 9965 68184
rect 2363 68153 2375 68156
rect 2317 68147 2375 68153
rect 3344 68116 3372 68156
rect 9953 68153 9965 68156
rect 9999 68153 10011 68187
rect 9953 68147 10011 68153
rect 2240 68088 3372 68116
rect 3421 68119 3479 68125
rect 3421 68085 3433 68119
rect 3467 68116 3479 68119
rect 8478 68116 8484 68128
rect 3467 68088 8484 68116
rect 3467 68085 3479 68088
rect 3421 68079 3479 68085
rect 8478 68076 8484 68088
rect 8536 68076 8542 68128
rect 1104 68026 10856 68048
rect 1104 67974 2582 68026
rect 2634 67974 2646 68026
rect 2698 67974 2710 68026
rect 2762 67974 2774 68026
rect 2826 67974 2838 68026
rect 2890 67974 5845 68026
rect 5897 67974 5909 68026
rect 5961 67974 5973 68026
rect 6025 67974 6037 68026
rect 6089 67974 6101 68026
rect 6153 67974 9109 68026
rect 9161 67974 9173 68026
rect 9225 67974 9237 68026
rect 9289 67974 9301 68026
rect 9353 67974 9365 68026
rect 9417 67974 10856 68026
rect 1104 67952 10856 67974
rect 845 67915 903 67921
rect 845 67881 857 67915
rect 891 67912 903 67915
rect 3786 67912 3792 67924
rect 891 67884 3792 67912
rect 891 67881 903 67884
rect 845 67875 903 67881
rect 3786 67872 3792 67884
rect 3844 67872 3850 67924
rect 937 67847 995 67853
rect 937 67813 949 67847
rect 983 67844 995 67847
rect 1394 67844 1400 67856
rect 983 67816 1400 67844
rect 983 67813 995 67816
rect 937 67807 995 67813
rect 1394 67804 1400 67816
rect 1452 67804 1458 67856
rect 3142 67804 3148 67856
rect 3200 67844 3206 67856
rect 3418 67844 3424 67856
rect 3200 67816 3424 67844
rect 3200 67804 3206 67816
rect 3418 67804 3424 67816
rect 3476 67804 3482 67856
rect 1394 67708 1400 67720
rect 1355 67680 1400 67708
rect 1394 67668 1400 67680
rect 1452 67668 1458 67720
rect 1673 67711 1731 67717
rect 1673 67677 1685 67711
rect 1719 67708 1731 67711
rect 1854 67708 1860 67720
rect 1719 67680 1860 67708
rect 1719 67677 1731 67680
rect 1673 67671 1731 67677
rect 1854 67668 1860 67680
rect 1912 67668 1918 67720
rect 10137 67711 10195 67717
rect 10137 67677 10149 67711
rect 10183 67677 10195 67711
rect 10137 67671 10195 67677
rect 2958 67640 2964 67652
rect 2919 67612 2964 67640
rect 2958 67600 2964 67612
rect 3016 67600 3022 67652
rect 3050 67600 3056 67652
rect 3108 67640 3114 67652
rect 3145 67643 3203 67649
rect 3145 67640 3157 67643
rect 3108 67612 3157 67640
rect 3108 67600 3114 67612
rect 3145 67609 3157 67612
rect 3191 67640 3203 67643
rect 3878 67640 3884 67652
rect 3191 67612 3884 67640
rect 3191 67609 3203 67612
rect 3145 67603 3203 67609
rect 3878 67600 3884 67612
rect 3936 67600 3942 67652
rect 10152 67584 10180 67671
rect 9950 67572 9956 67584
rect 9911 67544 9956 67572
rect 9950 67532 9956 67544
rect 10008 67532 10014 67584
rect 10134 67532 10140 67584
rect 10192 67532 10198 67584
rect 1104 67482 10856 67504
rect 1104 67430 4213 67482
rect 4265 67430 4277 67482
rect 4329 67430 4341 67482
rect 4393 67430 4405 67482
rect 4457 67430 4469 67482
rect 4521 67430 7477 67482
rect 7529 67430 7541 67482
rect 7593 67430 7605 67482
rect 7657 67430 7669 67482
rect 7721 67430 7733 67482
rect 7785 67430 10856 67482
rect 1104 67408 10856 67430
rect 2961 67371 3019 67377
rect 2961 67337 2973 67371
rect 3007 67368 3019 67371
rect 3326 67368 3332 67380
rect 3007 67340 3332 67368
rect 3007 67337 3019 67340
rect 2961 67331 3019 67337
rect 3326 67328 3332 67340
rect 3384 67328 3390 67380
rect 2133 67303 2191 67309
rect 2133 67269 2145 67303
rect 2179 67300 2191 67303
rect 9950 67300 9956 67312
rect 2179 67272 9956 67300
rect 2179 67269 2191 67272
rect 2133 67263 2191 67269
rect 9950 67260 9956 67272
rect 10008 67260 10014 67312
rect 1486 67192 1492 67244
rect 1544 67232 1550 67244
rect 1989 67235 2047 67241
rect 1989 67232 2001 67235
rect 1544 67204 2001 67232
rect 1544 67192 1550 67204
rect 1989 67201 2001 67204
rect 2035 67201 2047 67235
rect 1989 67195 2047 67201
rect 2225 67235 2283 67241
rect 2225 67201 2237 67235
rect 2271 67232 2283 67235
rect 2314 67232 2320 67244
rect 2271 67204 2320 67232
rect 2271 67201 2283 67204
rect 2225 67195 2283 67201
rect 2314 67192 2320 67204
rect 2372 67192 2378 67244
rect 2409 67235 2467 67241
rect 2409 67201 2421 67235
rect 2455 67201 2467 67235
rect 2409 67195 2467 67201
rect 1670 67124 1676 67176
rect 1728 67164 1734 67176
rect 2424 67164 2452 67195
rect 2958 67192 2964 67244
rect 3016 67232 3022 67244
rect 3053 67235 3111 67241
rect 3053 67232 3065 67235
rect 3016 67204 3065 67232
rect 3016 67192 3022 67204
rect 3053 67201 3065 67204
rect 3099 67232 3111 67235
rect 3142 67232 3148 67244
rect 3099 67204 3148 67232
rect 3099 67201 3111 67204
rect 3053 67195 3111 67201
rect 3142 67192 3148 67204
rect 3200 67192 3206 67244
rect 1728 67136 2452 67164
rect 1728 67124 1734 67136
rect 1857 67099 1915 67105
rect 1857 67065 1869 67099
rect 1903 67096 1915 67099
rect 5350 67096 5356 67108
rect 1903 67068 5356 67096
rect 1903 67065 1915 67068
rect 1857 67059 1915 67065
rect 5350 67056 5356 67068
rect 5408 67056 5414 67108
rect 1104 66938 10856 66960
rect 1104 66886 2582 66938
rect 2634 66886 2646 66938
rect 2698 66886 2710 66938
rect 2762 66886 2774 66938
rect 2826 66886 2838 66938
rect 2890 66886 5845 66938
rect 5897 66886 5909 66938
rect 5961 66886 5973 66938
rect 6025 66886 6037 66938
rect 6089 66886 6101 66938
rect 6153 66886 9109 66938
rect 9161 66886 9173 66938
rect 9225 66886 9237 66938
rect 9289 66886 9301 66938
rect 9353 66886 9365 66938
rect 9417 66886 10856 66938
rect 1104 66864 10856 66886
rect 1673 66623 1731 66629
rect 1673 66589 1685 66623
rect 1719 66589 1731 66623
rect 2314 66620 2320 66632
rect 2275 66592 2320 66620
rect 1673 66583 1731 66589
rect 1688 66552 1716 66583
rect 2314 66580 2320 66592
rect 2372 66580 2378 66632
rect 2958 66620 2964 66632
rect 2919 66592 2964 66620
rect 2958 66580 2964 66592
rect 3016 66580 3022 66632
rect 3326 66580 3332 66632
rect 3384 66620 3390 66632
rect 3602 66620 3608 66632
rect 3384 66592 3608 66620
rect 3384 66580 3390 66592
rect 3602 66580 3608 66592
rect 3660 66580 3666 66632
rect 10134 66620 10140 66632
rect 10095 66592 10140 66620
rect 10134 66580 10140 66592
rect 10192 66580 10198 66632
rect 6914 66552 6920 66564
rect 1688 66524 6920 66552
rect 6914 66512 6920 66524
rect 6972 66512 6978 66564
rect 1486 66484 1492 66496
rect 1447 66456 1492 66484
rect 1486 66444 1492 66456
rect 1544 66444 1550 66496
rect 2130 66484 2136 66496
rect 2091 66456 2136 66484
rect 2130 66444 2136 66456
rect 2188 66444 2194 66496
rect 2777 66487 2835 66493
rect 2777 66453 2789 66487
rect 2823 66484 2835 66487
rect 3602 66484 3608 66496
rect 2823 66456 3608 66484
rect 2823 66453 2835 66456
rect 2777 66447 2835 66453
rect 3602 66444 3608 66456
rect 3660 66444 3666 66496
rect 9950 66484 9956 66496
rect 9911 66456 9956 66484
rect 9950 66444 9956 66456
rect 10008 66444 10014 66496
rect 1104 66394 10856 66416
rect 1104 66342 4213 66394
rect 4265 66342 4277 66394
rect 4329 66342 4341 66394
rect 4393 66342 4405 66394
rect 4457 66342 4469 66394
rect 4521 66342 7477 66394
rect 7529 66342 7541 66394
rect 7593 66342 7605 66394
rect 7657 66342 7669 66394
rect 7721 66342 7733 66394
rect 7785 66342 10856 66394
rect 1104 66320 10856 66342
rect 753 66147 811 66153
rect 753 66113 765 66147
rect 799 66144 811 66147
rect 1673 66147 1731 66153
rect 1673 66144 1685 66147
rect 799 66116 1685 66144
rect 799 66113 811 66116
rect 753 66107 811 66113
rect 1673 66113 1685 66116
rect 1719 66113 1731 66147
rect 10134 66144 10140 66156
rect 10095 66116 10140 66144
rect 1673 66107 1731 66113
rect 10134 66104 10140 66116
rect 10192 66104 10198 66156
rect 1394 66076 1400 66088
rect 1355 66048 1400 66076
rect 1394 66036 1400 66048
rect 1452 66036 1458 66088
rect 9858 65900 9864 65952
rect 9916 65940 9922 65952
rect 9953 65943 10011 65949
rect 9953 65940 9965 65943
rect 9916 65912 9965 65940
rect 9916 65900 9922 65912
rect 9953 65909 9965 65912
rect 9999 65909 10011 65943
rect 9953 65903 10011 65909
rect 1104 65850 10856 65872
rect 1104 65798 2582 65850
rect 2634 65798 2646 65850
rect 2698 65798 2710 65850
rect 2762 65798 2774 65850
rect 2826 65798 2838 65850
rect 2890 65798 5845 65850
rect 5897 65798 5909 65850
rect 5961 65798 5973 65850
rect 6025 65798 6037 65850
rect 6089 65798 6101 65850
rect 6153 65798 9109 65850
rect 9161 65798 9173 65850
rect 9225 65798 9237 65850
rect 9289 65798 9301 65850
rect 9353 65798 9365 65850
rect 9417 65798 10856 65850
rect 1104 65776 10856 65798
rect 1026 65492 1032 65544
rect 1084 65532 1090 65544
rect 1673 65535 1731 65541
rect 1673 65532 1685 65535
rect 1084 65504 1685 65532
rect 1084 65492 1090 65504
rect 1673 65501 1685 65504
rect 1719 65501 1731 65535
rect 1673 65495 1731 65501
rect 2133 65535 2191 65541
rect 2133 65501 2145 65535
rect 2179 65501 2191 65535
rect 2133 65495 2191 65501
rect 2869 65535 2927 65541
rect 2869 65501 2881 65535
rect 2915 65532 2927 65535
rect 5626 65532 5632 65544
rect 2915 65504 5632 65532
rect 2915 65501 2927 65504
rect 2869 65495 2927 65501
rect 474 65424 480 65476
rect 532 65464 538 65476
rect 2148 65464 2176 65495
rect 5626 65492 5632 65504
rect 5684 65492 5690 65544
rect 10134 65532 10140 65544
rect 10095 65504 10140 65532
rect 10134 65492 10140 65504
rect 10192 65492 10198 65544
rect 532 65436 2176 65464
rect 532 65424 538 65436
rect 1486 65396 1492 65408
rect 1447 65368 1492 65396
rect 1486 65356 1492 65368
rect 1544 65356 1550 65408
rect 2314 65396 2320 65408
rect 2275 65368 2320 65396
rect 2314 65356 2320 65368
rect 2372 65356 2378 65408
rect 3050 65396 3056 65408
rect 3011 65368 3056 65396
rect 3050 65356 3056 65368
rect 3108 65356 3114 65408
rect 9766 65356 9772 65408
rect 9824 65396 9830 65408
rect 9953 65399 10011 65405
rect 9953 65396 9965 65399
rect 9824 65368 9965 65396
rect 9824 65356 9830 65368
rect 9953 65365 9965 65368
rect 9999 65365 10011 65399
rect 9953 65359 10011 65365
rect 1104 65306 10856 65328
rect 1104 65254 4213 65306
rect 4265 65254 4277 65306
rect 4329 65254 4341 65306
rect 4393 65254 4405 65306
rect 4457 65254 4469 65306
rect 4521 65254 7477 65306
rect 7529 65254 7541 65306
rect 7593 65254 7605 65306
rect 7657 65254 7669 65306
rect 7721 65254 7733 65306
rect 7785 65254 10856 65306
rect 1104 65232 10856 65254
rect 1946 65124 1952 65136
rect 1907 65096 1952 65124
rect 1946 65084 1952 65096
rect 2004 65084 2010 65136
rect 2041 65127 2099 65133
rect 2041 65093 2053 65127
rect 2087 65124 2099 65127
rect 9950 65124 9956 65136
rect 2087 65096 9956 65124
rect 2087 65093 2099 65096
rect 2041 65087 2099 65093
rect 9950 65084 9956 65096
rect 10008 65084 10014 65136
rect 1670 65016 1676 65068
rect 1728 65056 1734 65068
rect 1765 65059 1823 65065
rect 1765 65056 1777 65059
rect 1728 65028 1777 65056
rect 1728 65016 1734 65028
rect 1765 65025 1777 65028
rect 1811 65025 1823 65059
rect 1765 65019 1823 65025
rect 2138 65059 2196 65065
rect 2138 65025 2150 65059
rect 2184 65025 2196 65059
rect 3145 65059 3203 65065
rect 3145 65056 3157 65059
rect 2138 65019 2196 65025
rect 2746 65028 3157 65056
rect 1394 64948 1400 65000
rect 1452 64988 1458 65000
rect 1946 64988 1952 65000
rect 1452 64960 1952 64988
rect 1452 64948 1458 64960
rect 1946 64948 1952 64960
rect 2004 64988 2010 65000
rect 2148 64988 2176 65019
rect 2746 64988 2774 65028
rect 3145 65025 3157 65028
rect 3191 65025 3203 65059
rect 3145 65019 3203 65025
rect 2004 64960 2774 64988
rect 2869 64991 2927 64997
rect 2004 64948 2010 64960
rect 2869 64957 2881 64991
rect 2915 64988 2927 64991
rect 3050 64988 3056 65000
rect 2915 64960 3056 64988
rect 2915 64957 2927 64960
rect 2869 64951 2927 64957
rect 3050 64948 3056 64960
rect 3108 64948 3114 65000
rect 2317 64923 2375 64929
rect 2317 64889 2329 64923
rect 2363 64920 2375 64923
rect 11333 64923 11391 64929
rect 11333 64920 11345 64923
rect 2363 64892 11345 64920
rect 2363 64889 2375 64892
rect 2317 64883 2375 64889
rect 11333 64889 11345 64892
rect 11379 64889 11391 64923
rect 11333 64883 11391 64889
rect 1104 64762 10856 64784
rect 1104 64710 2582 64762
rect 2634 64710 2646 64762
rect 2698 64710 2710 64762
rect 2762 64710 2774 64762
rect 2826 64710 2838 64762
rect 2890 64710 5845 64762
rect 5897 64710 5909 64762
rect 5961 64710 5973 64762
rect 6025 64710 6037 64762
rect 6089 64710 6101 64762
rect 6153 64710 9109 64762
rect 9161 64710 9173 64762
rect 9225 64710 9237 64762
rect 9289 64710 9301 64762
rect 9353 64710 9365 64762
rect 9417 64710 10856 64762
rect 1104 64688 10856 64710
rect 1670 64540 1676 64592
rect 1728 64540 1734 64592
rect 1688 64512 1716 64540
rect 2406 64512 2412 64524
rect 1688 64484 2412 64512
rect 2406 64472 2412 64484
rect 2464 64512 2470 64524
rect 2593 64515 2651 64521
rect 2593 64512 2605 64515
rect 2464 64484 2605 64512
rect 2464 64472 2470 64484
rect 2593 64481 2605 64484
rect 2639 64481 2651 64515
rect 2593 64475 2651 64481
rect 9861 64515 9919 64521
rect 9861 64481 9873 64515
rect 9907 64512 9919 64515
rect 11425 64515 11483 64521
rect 11425 64512 11437 64515
rect 9907 64484 11437 64512
rect 9907 64481 9919 64484
rect 9861 64475 9919 64481
rect 11425 64481 11437 64484
rect 11471 64481 11483 64515
rect 11425 64475 11483 64481
rect 1673 64447 1731 64453
rect 1673 64413 1685 64447
rect 1719 64413 1731 64447
rect 1673 64407 1731 64413
rect 2317 64447 2375 64453
rect 2317 64413 2329 64447
rect 2363 64413 2375 64447
rect 10134 64444 10140 64456
rect 10095 64416 10140 64444
rect 2317 64407 2375 64413
rect 1394 64268 1400 64320
rect 1452 64308 1458 64320
rect 1489 64311 1547 64317
rect 1489 64308 1501 64311
rect 1452 64280 1501 64308
rect 1452 64268 1458 64280
rect 1489 64277 1501 64280
rect 1535 64277 1547 64311
rect 1688 64308 1716 64407
rect 2332 64376 2360 64407
rect 10134 64404 10140 64416
rect 10192 64404 10198 64456
rect 3418 64376 3424 64388
rect 2332 64348 3424 64376
rect 3418 64336 3424 64348
rect 3476 64336 3482 64388
rect 3786 64308 3792 64320
rect 1688 64280 3792 64308
rect 1489 64271 1547 64277
rect 3786 64268 3792 64280
rect 3844 64268 3850 64320
rect 1104 64218 10856 64240
rect 1104 64166 4213 64218
rect 4265 64166 4277 64218
rect 4329 64166 4341 64218
rect 4393 64166 4405 64218
rect 4457 64166 4469 64218
rect 4521 64166 7477 64218
rect 7529 64166 7541 64218
rect 7593 64166 7605 64218
rect 7657 64166 7669 64218
rect 7721 64166 7733 64218
rect 7785 64166 10856 64218
rect 1104 64144 10856 64166
rect 9858 64104 9864 64116
rect 2746 64076 9864 64104
rect 2225 64039 2283 64045
rect 2225 64005 2237 64039
rect 2271 64036 2283 64039
rect 2746 64036 2774 64076
rect 9858 64064 9864 64076
rect 9916 64064 9922 64116
rect 2271 64008 2774 64036
rect 2271 64005 2283 64008
rect 2225 63999 2283 64005
rect 1946 63928 1952 63980
rect 2004 63968 2010 63980
rect 2081 63971 2139 63977
rect 2081 63968 2093 63971
rect 2004 63940 2093 63968
rect 2004 63928 2010 63940
rect 2081 63937 2093 63940
rect 2127 63937 2139 63971
rect 2081 63931 2139 63937
rect 2317 63971 2375 63977
rect 2317 63937 2329 63971
rect 2363 63937 2375 63971
rect 2317 63931 2375 63937
rect 1578 63860 1584 63912
rect 1636 63900 1642 63912
rect 2332 63900 2360 63931
rect 2406 63928 2412 63980
rect 2464 63968 2470 63980
rect 2501 63971 2559 63977
rect 2501 63968 2513 63971
rect 2464 63940 2513 63968
rect 2464 63928 2470 63940
rect 2501 63937 2513 63940
rect 2547 63937 2559 63971
rect 2501 63931 2559 63937
rect 2961 63971 3019 63977
rect 2961 63937 2973 63971
rect 3007 63937 3019 63971
rect 2961 63931 3019 63937
rect 3697 63971 3755 63977
rect 3697 63937 3709 63971
rect 3743 63968 3755 63971
rect 5074 63968 5080 63980
rect 3743 63940 5080 63968
rect 3743 63937 3755 63940
rect 3697 63931 3755 63937
rect 1636 63872 2360 63900
rect 2976 63900 3004 63931
rect 5074 63928 5080 63940
rect 5132 63928 5138 63980
rect 9861 63971 9919 63977
rect 9861 63937 9873 63971
rect 9907 63968 9919 63971
rect 11241 63971 11299 63977
rect 11241 63968 11253 63971
rect 9907 63940 11253 63968
rect 9907 63937 9919 63940
rect 9861 63931 9919 63937
rect 11241 63937 11253 63940
rect 11287 63937 11299 63971
rect 11241 63931 11299 63937
rect 5166 63900 5172 63912
rect 2976 63872 5172 63900
rect 1636 63860 1642 63872
rect 5166 63860 5172 63872
rect 5224 63860 5230 63912
rect 10134 63900 10140 63912
rect 10095 63872 10140 63900
rect 10134 63860 10140 63872
rect 10192 63860 10198 63912
rect 3878 63832 3884 63844
rect 2746 63804 3280 63832
rect 3839 63804 3884 63832
rect 1949 63767 2007 63773
rect 1949 63733 1961 63767
rect 1995 63764 2007 63767
rect 2746 63764 2774 63804
rect 3142 63764 3148 63776
rect 1995 63736 2774 63764
rect 3103 63736 3148 63764
rect 1995 63733 2007 63736
rect 1949 63727 2007 63733
rect 3142 63724 3148 63736
rect 3200 63724 3206 63776
rect 3252 63764 3280 63804
rect 3878 63792 3884 63804
rect 3936 63792 3942 63844
rect 6270 63764 6276 63776
rect 3252 63736 6276 63764
rect 6270 63724 6276 63736
rect 6328 63724 6334 63776
rect 1104 63674 10856 63696
rect 1104 63622 2582 63674
rect 2634 63622 2646 63674
rect 2698 63622 2710 63674
rect 2762 63622 2774 63674
rect 2826 63622 2838 63674
rect 2890 63622 5845 63674
rect 5897 63622 5909 63674
rect 5961 63622 5973 63674
rect 6025 63622 6037 63674
rect 6089 63622 6101 63674
rect 6153 63622 9109 63674
rect 9161 63622 9173 63674
rect 9225 63622 9237 63674
rect 9289 63622 9301 63674
rect 9353 63622 9365 63674
rect 9417 63622 10856 63674
rect 1104 63600 10856 63622
rect 1949 63563 2007 63569
rect 1949 63529 1961 63563
rect 1995 63560 2007 63563
rect 5442 63560 5448 63572
rect 1995 63532 5448 63560
rect 1995 63529 2007 63532
rect 1949 63523 2007 63529
rect 5442 63520 5448 63532
rect 5500 63520 5506 63572
rect 2593 63495 2651 63501
rect 2593 63461 2605 63495
rect 2639 63492 2651 63495
rect 8570 63492 8576 63504
rect 2639 63464 8576 63492
rect 2639 63461 2651 63464
rect 2593 63455 2651 63461
rect 8570 63452 8576 63464
rect 8628 63452 8634 63504
rect 1670 63424 1676 63436
rect 1412 63396 1676 63424
rect 1412 63365 1440 63396
rect 1670 63384 1676 63396
rect 1728 63384 1734 63436
rect 2866 63384 2872 63436
rect 2924 63384 2930 63436
rect 1397 63359 1455 63365
rect 1397 63325 1409 63359
rect 1443 63325 1455 63359
rect 1397 63319 1455 63325
rect 1817 63359 1875 63365
rect 1817 63325 1829 63359
rect 1863 63356 1875 63359
rect 1946 63356 1952 63368
rect 1863 63328 1952 63356
rect 1863 63325 1875 63328
rect 1817 63319 1875 63325
rect 1946 63316 1952 63328
rect 2004 63316 2010 63368
rect 2406 63316 2412 63368
rect 2464 63356 2470 63368
rect 2725 63359 2783 63365
rect 2725 63356 2737 63359
rect 2464 63328 2737 63356
rect 2464 63316 2470 63328
rect 2725 63325 2737 63328
rect 2771 63325 2783 63359
rect 2884 63356 2912 63384
rect 3007 63359 3065 63365
rect 3007 63356 3019 63359
rect 2884 63328 3019 63356
rect 2725 63319 2783 63325
rect 3007 63325 3019 63328
rect 3053 63325 3065 63359
rect 3007 63319 3065 63325
rect 3099 63359 3157 63365
rect 3099 63325 3111 63359
rect 3145 63356 3157 63359
rect 3789 63359 3847 63365
rect 3145 63328 3372 63356
rect 3145 63325 3157 63328
rect 3099 63319 3157 63325
rect 1581 63291 1639 63297
rect 1581 63257 1593 63291
rect 1627 63257 1639 63291
rect 1581 63251 1639 63257
rect 1596 63220 1624 63251
rect 1670 63248 1676 63300
rect 1728 63288 1734 63300
rect 2866 63288 2872 63300
rect 1728 63260 1773 63288
rect 2827 63260 2872 63288
rect 1728 63248 1734 63260
rect 2866 63248 2872 63260
rect 2924 63248 2930 63300
rect 3344 63288 3372 63328
rect 3789 63325 3801 63359
rect 3835 63356 3847 63359
rect 5718 63356 5724 63368
rect 3835 63328 5724 63356
rect 3835 63325 3847 63328
rect 3789 63319 3847 63325
rect 5718 63316 5724 63328
rect 5776 63316 5782 63368
rect 3878 63288 3884 63300
rect 3344 63260 3884 63288
rect 3878 63248 3884 63260
rect 3936 63248 3942 63300
rect 4062 63248 4068 63300
rect 4120 63288 4126 63300
rect 9950 63288 9956 63300
rect 4120 63260 9956 63288
rect 4120 63248 4126 63260
rect 9950 63248 9956 63260
rect 10008 63248 10014 63300
rect 2314 63220 2320 63232
rect 1596 63192 2320 63220
rect 2314 63180 2320 63192
rect 2372 63180 2378 63232
rect 3970 63220 3976 63232
rect 3931 63192 3976 63220
rect 3970 63180 3976 63192
rect 4028 63180 4034 63232
rect 1104 63130 10856 63152
rect 1104 63078 4213 63130
rect 4265 63078 4277 63130
rect 4329 63078 4341 63130
rect 4393 63078 4405 63130
rect 4457 63078 4469 63130
rect 4521 63078 7477 63130
rect 7529 63078 7541 63130
rect 7593 63078 7605 63130
rect 7657 63078 7669 63130
rect 7721 63078 7733 63130
rect 7785 63078 10856 63130
rect 1104 63056 10856 63078
rect 1670 62976 1676 63028
rect 1728 63016 1734 63028
rect 9950 63016 9956 63028
rect 1728 62988 2912 63016
rect 9911 62988 9956 63016
rect 1728 62976 1734 62988
rect 2314 62908 2320 62960
rect 2372 62948 2378 62960
rect 2884 62948 2912 62988
rect 9950 62976 9956 62988
rect 10008 62976 10014 63028
rect 9766 62948 9772 62960
rect 2372 62920 2820 62948
rect 2884 62920 9772 62948
rect 2372 62908 2378 62920
rect 1578 62840 1584 62892
rect 1636 62880 1642 62892
rect 1673 62883 1731 62889
rect 1673 62880 1685 62883
rect 1636 62852 1685 62880
rect 1636 62840 1642 62852
rect 1673 62849 1685 62852
rect 1719 62849 1731 62883
rect 1673 62843 1731 62849
rect 2409 62883 2467 62889
rect 2409 62849 2421 62883
rect 2455 62849 2467 62883
rect 2792 62880 2820 62920
rect 9766 62908 9772 62920
rect 9824 62908 9830 62960
rect 3145 62883 3203 62889
rect 3145 62880 3157 62883
rect 2792 62852 3157 62880
rect 2409 62843 2467 62849
rect 3145 62849 3157 62852
rect 3191 62849 3203 62883
rect 3145 62843 3203 62849
rect 4157 62883 4215 62889
rect 4157 62849 4169 62883
rect 4203 62880 4215 62883
rect 4982 62880 4988 62892
rect 4203 62852 4988 62880
rect 4203 62849 4215 62852
rect 4157 62843 4215 62849
rect 934 62772 940 62824
rect 992 62812 998 62824
rect 2314 62812 2320 62824
rect 992 62784 2320 62812
rect 992 62772 998 62784
rect 2314 62772 2320 62784
rect 2372 62772 2378 62824
rect 1486 62676 1492 62688
rect 1447 62648 1492 62676
rect 1486 62636 1492 62648
rect 1544 62636 1550 62688
rect 2222 62676 2228 62688
rect 2183 62648 2228 62676
rect 2222 62636 2228 62648
rect 2280 62636 2286 62688
rect 2424 62676 2452 62843
rect 4982 62840 4988 62852
rect 5040 62840 5046 62892
rect 10134 62880 10140 62892
rect 10095 62852 10140 62880
rect 10134 62840 10140 62852
rect 10192 62840 10198 62892
rect 2869 62815 2927 62821
rect 2869 62781 2881 62815
rect 2915 62812 2927 62815
rect 3050 62812 3056 62824
rect 2915 62784 3056 62812
rect 2915 62781 2927 62784
rect 2869 62775 2927 62781
rect 3050 62772 3056 62784
rect 3108 62812 3114 62824
rect 4249 62815 4307 62821
rect 4249 62812 4261 62815
rect 3108 62784 4261 62812
rect 3108 62772 3114 62784
rect 4249 62781 4261 62784
rect 4295 62781 4307 62815
rect 4249 62775 4307 62781
rect 5442 62704 5448 62756
rect 5500 62744 5506 62756
rect 11609 62747 11667 62753
rect 11609 62744 11621 62747
rect 5500 62716 11621 62744
rect 5500 62704 5506 62716
rect 11609 62713 11621 62716
rect 11655 62713 11667 62747
rect 11609 62707 11667 62713
rect 3050 62676 3056 62688
rect 2424 62648 3056 62676
rect 3050 62636 3056 62648
rect 3108 62636 3114 62688
rect 1104 62586 10856 62608
rect 1104 62534 2582 62586
rect 2634 62534 2646 62586
rect 2698 62534 2710 62586
rect 2762 62534 2774 62586
rect 2826 62534 2838 62586
rect 2890 62534 5845 62586
rect 5897 62534 5909 62586
rect 5961 62534 5973 62586
rect 6025 62534 6037 62586
rect 6089 62534 6101 62586
rect 6153 62534 9109 62586
rect 9161 62534 9173 62586
rect 9225 62534 9237 62586
rect 9289 62534 9301 62586
rect 9353 62534 9365 62586
rect 9417 62534 10856 62586
rect 1104 62512 10856 62534
rect 658 62432 664 62484
rect 716 62472 722 62484
rect 1949 62475 2007 62481
rect 1949 62472 1961 62475
rect 716 62444 1961 62472
rect 716 62432 722 62444
rect 1949 62441 1961 62444
rect 1995 62441 2007 62475
rect 1949 62435 2007 62441
rect 2593 62475 2651 62481
rect 2593 62441 2605 62475
rect 2639 62472 2651 62475
rect 5442 62472 5448 62484
rect 2639 62444 5448 62472
rect 2639 62441 2651 62444
rect 2593 62435 2651 62441
rect 5442 62432 5448 62444
rect 5500 62432 5506 62484
rect 1394 62364 1400 62416
rect 1452 62404 1458 62416
rect 1762 62404 1768 62416
rect 1452 62376 1768 62404
rect 1452 62364 1458 62376
rect 1762 62364 1768 62376
rect 1820 62364 1826 62416
rect 937 62339 995 62345
rect 937 62305 949 62339
rect 983 62336 995 62339
rect 9674 62336 9680 62348
rect 983 62308 1624 62336
rect 983 62305 995 62308
rect 937 62299 995 62305
rect 1596 62277 1624 62308
rect 1688 62308 9680 62336
rect 1688 62277 1716 62308
rect 9674 62296 9680 62308
rect 9732 62296 9738 62348
rect 1397 62271 1455 62277
rect 1397 62237 1409 62271
rect 1443 62237 1455 62271
rect 1397 62231 1455 62237
rect 1581 62271 1639 62277
rect 1581 62237 1593 62271
rect 1627 62237 1639 62271
rect 1581 62231 1639 62237
rect 1673 62271 1731 62277
rect 1673 62237 1685 62271
rect 1719 62237 1731 62271
rect 1673 62231 1731 62237
rect 1412 62132 1440 62231
rect 1762 62228 1768 62280
rect 1820 62277 1826 62280
rect 1820 62268 1828 62277
rect 1820 62240 1865 62268
rect 1820 62231 1828 62240
rect 1820 62228 1826 62231
rect 2406 62228 2412 62280
rect 2464 62268 2470 62280
rect 2725 62271 2783 62277
rect 2725 62268 2737 62271
rect 2464 62240 2737 62268
rect 2464 62228 2470 62240
rect 2725 62237 2737 62240
rect 2771 62237 2783 62271
rect 2725 62231 2783 62237
rect 3145 62271 3203 62277
rect 3145 62237 3157 62271
rect 3191 62268 3203 62271
rect 3878 62268 3884 62280
rect 3191 62240 3884 62268
rect 3191 62237 3203 62240
rect 3145 62231 3203 62237
rect 3878 62228 3884 62240
rect 3936 62228 3942 62280
rect 10134 62268 10140 62280
rect 10095 62240 10140 62268
rect 10134 62228 10140 62240
rect 10192 62228 10198 62280
rect 2869 62203 2927 62209
rect 2869 62169 2881 62203
rect 2915 62169 2927 62203
rect 2869 62163 2927 62169
rect 2961 62203 3019 62209
rect 2961 62169 2973 62203
rect 3007 62200 3019 62203
rect 3510 62200 3516 62212
rect 3007 62172 3516 62200
rect 3007 62169 3019 62172
rect 2961 62163 3019 62169
rect 1946 62132 1952 62144
rect 1412 62104 1952 62132
rect 1946 62092 1952 62104
rect 2004 62092 2010 62144
rect 2884 62132 2912 62163
rect 3510 62160 3516 62172
rect 3568 62160 3574 62212
rect 9953 62135 10011 62141
rect 9953 62132 9965 62135
rect 2884 62104 9965 62132
rect 9953 62101 9965 62104
rect 9999 62101 10011 62135
rect 9953 62095 10011 62101
rect 1104 62042 10856 62064
rect 1104 61990 4213 62042
rect 4265 61990 4277 62042
rect 4329 61990 4341 62042
rect 4393 61990 4405 62042
rect 4457 61990 4469 62042
rect 4521 61990 7477 62042
rect 7529 61990 7541 62042
rect 7593 61990 7605 62042
rect 7657 61990 7669 62042
rect 7721 61990 7733 62042
rect 7785 61990 10856 62042
rect 1104 61968 10856 61990
rect 1966 61931 2024 61937
rect 1966 61897 1978 61931
rect 2012 61928 2024 61931
rect 4062 61928 4068 61940
rect 2012 61900 4068 61928
rect 2012 61897 2024 61900
rect 1966 61891 2024 61897
rect 4062 61888 4068 61900
rect 4120 61888 4126 61940
rect 2958 61820 2964 61872
rect 3016 61860 3022 61872
rect 3142 61860 3148 61872
rect 3016 61832 3148 61860
rect 3016 61820 3022 61832
rect 3142 61820 3148 61832
rect 3200 61820 3206 61872
rect 1397 61795 1455 61801
rect 1397 61761 1409 61795
rect 1443 61792 1455 61795
rect 1581 61795 1639 61801
rect 1443 61764 1532 61792
rect 1443 61761 1455 61764
rect 1397 61755 1455 61761
rect 1504 61588 1532 61764
rect 1581 61761 1593 61795
rect 1627 61761 1639 61795
rect 1581 61755 1639 61761
rect 1673 61795 1731 61801
rect 1673 61761 1685 61795
rect 1719 61761 1731 61795
rect 1673 61755 1731 61761
rect 1596 61656 1624 61755
rect 1688 61724 1716 61755
rect 1762 61752 1768 61804
rect 1820 61801 1826 61804
rect 1820 61792 1828 61801
rect 1820 61764 1865 61792
rect 1820 61755 1828 61764
rect 1820 61752 1826 61755
rect 2038 61752 2044 61804
rect 2096 61792 2102 61804
rect 2501 61795 2559 61801
rect 2501 61792 2513 61795
rect 2096 61764 2513 61792
rect 2096 61752 2102 61764
rect 2501 61761 2513 61764
rect 2547 61761 2559 61795
rect 10134 61792 10140 61804
rect 10095 61764 10140 61792
rect 2501 61755 2559 61761
rect 10134 61752 10140 61764
rect 10192 61752 10198 61804
rect 9766 61724 9772 61736
rect 1688 61696 9772 61724
rect 9766 61684 9772 61696
rect 9824 61684 9830 61736
rect 3694 61656 3700 61668
rect 1596 61628 3700 61656
rect 3694 61616 3700 61628
rect 3752 61616 3758 61668
rect 1946 61588 1952 61600
rect 1504 61560 1952 61588
rect 1946 61548 1952 61560
rect 2004 61548 2010 61600
rect 2685 61591 2743 61597
rect 2685 61557 2697 61591
rect 2731 61588 2743 61591
rect 2958 61588 2964 61600
rect 2731 61560 2964 61588
rect 2731 61557 2743 61560
rect 2685 61551 2743 61557
rect 2958 61548 2964 61560
rect 3016 61548 3022 61600
rect 9950 61588 9956 61600
rect 9911 61560 9956 61588
rect 9950 61548 9956 61560
rect 10008 61548 10014 61600
rect 1104 61498 10856 61520
rect 1104 61446 2582 61498
rect 2634 61446 2646 61498
rect 2698 61446 2710 61498
rect 2762 61446 2774 61498
rect 2826 61446 2838 61498
rect 2890 61446 5845 61498
rect 5897 61446 5909 61498
rect 5961 61446 5973 61498
rect 6025 61446 6037 61498
rect 6089 61446 6101 61498
rect 6153 61446 9109 61498
rect 9161 61446 9173 61498
rect 9225 61446 9237 61498
rect 9289 61446 9301 61498
rect 9353 61446 9365 61498
rect 9417 61446 10856 61498
rect 1104 61424 10856 61446
rect 1762 61344 1768 61396
rect 1820 61384 1826 61396
rect 2130 61384 2136 61396
rect 1820 61356 2136 61384
rect 1820 61344 1826 61356
rect 2130 61344 2136 61356
rect 2188 61344 2194 61396
rect 1489 61319 1547 61325
rect 1489 61285 1501 61319
rect 1535 61316 1547 61319
rect 11517 61319 11575 61325
rect 11517 61316 11529 61319
rect 1535 61288 11529 61316
rect 1535 61285 1547 61288
rect 1489 61279 1547 61285
rect 11517 61285 11529 61288
rect 11563 61285 11575 61319
rect 11517 61279 11575 61285
rect 1946 61208 1952 61260
rect 2004 61248 2010 61260
rect 2004 61220 2084 61248
rect 2004 61208 2010 61220
rect 1670 61189 1676 61192
rect 1668 61180 1676 61189
rect 1631 61152 1676 61180
rect 1668 61143 1676 61152
rect 1670 61140 1676 61143
rect 1728 61140 1734 61192
rect 2056 61189 2084 61220
rect 1765 61183 1823 61189
rect 1765 61149 1777 61183
rect 1811 61180 1823 61183
rect 2041 61183 2099 61189
rect 1811 61152 1992 61180
rect 1811 61149 1823 61152
rect 1765 61143 1823 61149
rect 845 61115 903 61121
rect 845 61081 857 61115
rect 891 61112 903 61115
rect 1857 61115 1915 61121
rect 1857 61112 1869 61115
rect 891 61084 1869 61112
rect 891 61081 903 61084
rect 845 61075 903 61081
rect 1857 61081 1869 61084
rect 1903 61081 1915 61115
rect 1964 61112 1992 61152
rect 2041 61149 2053 61183
rect 2087 61149 2099 61183
rect 2041 61143 2099 61149
rect 2222 61140 2228 61192
rect 2280 61180 2286 61192
rect 2501 61183 2559 61189
rect 2501 61180 2513 61183
rect 2280 61152 2513 61180
rect 2280 61140 2286 61152
rect 2501 61149 2513 61152
rect 2547 61149 2559 61183
rect 2501 61143 2559 61149
rect 3418 61140 3424 61192
rect 3476 61180 3482 61192
rect 3789 61183 3847 61189
rect 3789 61180 3801 61183
rect 3476 61152 3801 61180
rect 3476 61140 3482 61152
rect 3789 61149 3801 61152
rect 3835 61149 3847 61183
rect 3789 61143 3847 61149
rect 9858 61112 9864 61124
rect 1964 61084 9864 61112
rect 1857 61075 1915 61081
rect 9858 61072 9864 61084
rect 9916 61072 9922 61124
rect 2685 61047 2743 61053
rect 2685 61013 2697 61047
rect 2731 61044 2743 61047
rect 2774 61044 2780 61056
rect 2731 61016 2780 61044
rect 2731 61013 2743 61016
rect 2685 61007 2743 61013
rect 2774 61004 2780 61016
rect 2832 61004 2838 61056
rect 3970 61044 3976 61056
rect 3931 61016 3976 61044
rect 3970 61004 3976 61016
rect 4028 61004 4034 61056
rect 1104 60954 10856 60976
rect 1104 60902 4213 60954
rect 4265 60902 4277 60954
rect 4329 60902 4341 60954
rect 4393 60902 4405 60954
rect 4457 60902 4469 60954
rect 4521 60902 7477 60954
rect 7529 60902 7541 60954
rect 7593 60902 7605 60954
rect 7657 60902 7669 60954
rect 7721 60902 7733 60954
rect 7785 60902 10856 60954
rect 1104 60880 10856 60902
rect 845 60843 903 60849
rect 845 60809 857 60843
rect 891 60840 903 60843
rect 1394 60840 1400 60852
rect 891 60812 1400 60840
rect 891 60809 903 60812
rect 845 60803 903 60809
rect 1394 60800 1400 60812
rect 1452 60800 1458 60852
rect 1854 60840 1860 60852
rect 1596 60812 1860 60840
rect 1596 60784 1624 60812
rect 1854 60800 1860 60812
rect 1912 60800 1918 60852
rect 2406 60800 2412 60852
rect 2464 60800 2470 60852
rect 3326 60840 3332 60852
rect 2516 60812 3332 60840
rect 1578 60732 1584 60784
rect 1636 60732 1642 60784
rect 2424 60772 2452 60800
rect 2516 60781 2544 60812
rect 3326 60800 3332 60812
rect 3384 60800 3390 60852
rect 2240 60744 2452 60772
rect 937 60707 995 60713
rect 937 60673 949 60707
rect 983 60704 995 60707
rect 1302 60704 1308 60716
rect 983 60676 1308 60704
rect 983 60673 995 60676
rect 937 60667 995 60673
rect 1302 60664 1308 60676
rect 1360 60664 1366 60716
rect 1673 60707 1731 60713
rect 1673 60673 1685 60707
rect 1719 60704 1731 60707
rect 1854 60704 1860 60716
rect 1719 60676 1860 60704
rect 1719 60673 1731 60676
rect 1673 60667 1731 60673
rect 1854 60664 1860 60676
rect 1912 60664 1918 60716
rect 1486 60500 1492 60512
rect 1447 60472 1492 60500
rect 1486 60460 1492 60472
rect 1544 60460 1550 60512
rect 2240 60500 2268 60744
rect 2317 60707 2375 60713
rect 2317 60673 2329 60707
rect 2363 60673 2375 60707
rect 2424 60704 2452 60744
rect 2501 60775 2559 60781
rect 2501 60741 2513 60775
rect 2547 60741 2559 60775
rect 2501 60735 2559 60741
rect 2593 60775 2651 60781
rect 2593 60741 2605 60775
rect 2639 60772 2651 60775
rect 9950 60772 9956 60784
rect 2639 60744 9956 60772
rect 2639 60741 2651 60744
rect 2593 60735 2651 60741
rect 9950 60732 9956 60744
rect 10008 60732 10014 60784
rect 2690 60707 2748 60713
rect 2690 60704 2702 60707
rect 2424 60676 2702 60704
rect 2317 60667 2375 60673
rect 2690 60673 2702 60676
rect 2736 60673 2748 60707
rect 2690 60667 2748 60673
rect 2332 60636 2360 60667
rect 3602 60664 3608 60716
rect 3660 60664 3666 60716
rect 10134 60704 10140 60716
rect 10095 60676 10140 60704
rect 10134 60664 10140 60676
rect 10192 60664 10198 60716
rect 3326 60636 3332 60648
rect 2332 60608 3332 60636
rect 3326 60596 3332 60608
rect 3384 60596 3390 60648
rect 3620 60512 3648 60664
rect 9766 60528 9772 60580
rect 9824 60568 9830 60580
rect 9953 60571 10011 60577
rect 9953 60568 9965 60571
rect 9824 60540 9965 60568
rect 9824 60528 9830 60540
rect 9953 60537 9965 60540
rect 9999 60537 10011 60571
rect 9953 60531 10011 60537
rect 2314 60500 2320 60512
rect 2240 60472 2320 60500
rect 2314 60460 2320 60472
rect 2372 60460 2378 60512
rect 2869 60503 2927 60509
rect 2869 60469 2881 60503
rect 2915 60500 2927 60503
rect 3510 60500 3516 60512
rect 2915 60472 3516 60500
rect 2915 60469 2927 60472
rect 2869 60463 2927 60469
rect 3510 60460 3516 60472
rect 3568 60460 3574 60512
rect 3602 60460 3608 60512
rect 3660 60460 3666 60512
rect 1104 60410 10856 60432
rect 1104 60358 2582 60410
rect 2634 60358 2646 60410
rect 2698 60358 2710 60410
rect 2762 60358 2774 60410
rect 2826 60358 2838 60410
rect 2890 60358 5845 60410
rect 5897 60358 5909 60410
rect 5961 60358 5973 60410
rect 6025 60358 6037 60410
rect 6089 60358 6101 60410
rect 6153 60358 9109 60410
rect 9161 60358 9173 60410
rect 9225 60358 9237 60410
rect 9289 60358 9301 60410
rect 9353 60358 9365 60410
rect 9417 60358 10856 60410
rect 1104 60336 10856 60358
rect 1854 60256 1860 60308
rect 1912 60296 1918 60308
rect 3970 60296 3976 60308
rect 1912 60268 3976 60296
rect 1912 60256 1918 60268
rect 3970 60256 3976 60268
rect 4028 60256 4034 60308
rect 9674 60256 9680 60308
rect 9732 60296 9738 60308
rect 9953 60299 10011 60305
rect 9953 60296 9965 60299
rect 9732 60268 9965 60296
rect 9732 60256 9738 60268
rect 9953 60265 9965 60268
rect 9999 60265 10011 60299
rect 9953 60259 10011 60265
rect 1670 60188 1676 60240
rect 1728 60228 1734 60240
rect 1728 60200 2544 60228
rect 1728 60188 1734 60200
rect 1964 60104 1992 60200
rect 2516 60169 2544 60200
rect 2501 60163 2559 60169
rect 2501 60129 2513 60163
rect 2547 60129 2559 60163
rect 2501 60123 2559 60129
rect 1673 60095 1731 60101
rect 1673 60061 1685 60095
rect 1719 60061 1731 60095
rect 1673 60055 1731 60061
rect 1302 59916 1308 59968
rect 1360 59956 1366 59968
rect 1489 59959 1547 59965
rect 1489 59956 1501 59959
rect 1360 59928 1501 59956
rect 1360 59916 1366 59928
rect 1489 59925 1501 59928
rect 1535 59925 1547 59959
rect 1688 59956 1716 60055
rect 1946 60052 1952 60104
rect 2004 60052 2010 60104
rect 2225 60095 2283 60101
rect 2225 60061 2237 60095
rect 2271 60061 2283 60095
rect 10134 60092 10140 60104
rect 10095 60064 10140 60092
rect 2225 60055 2283 60061
rect 2240 60024 2268 60055
rect 10134 60052 10140 60064
rect 10192 60052 10198 60104
rect 2958 60024 2964 60036
rect 2240 59996 2964 60024
rect 2958 59984 2964 59996
rect 3016 60024 3022 60036
rect 3142 60024 3148 60036
rect 3016 59996 3148 60024
rect 3016 59984 3022 59996
rect 3142 59984 3148 59996
rect 3200 59984 3206 60036
rect 2866 59956 2872 59968
rect 1688 59928 2872 59956
rect 1489 59919 1547 59925
rect 2866 59916 2872 59928
rect 2924 59916 2930 59968
rect 1104 59866 10856 59888
rect 1104 59814 4213 59866
rect 4265 59814 4277 59866
rect 4329 59814 4341 59866
rect 4393 59814 4405 59866
rect 4457 59814 4469 59866
rect 4521 59814 7477 59866
rect 7529 59814 7541 59866
rect 7593 59814 7605 59866
rect 7657 59814 7669 59866
rect 7721 59814 7733 59866
rect 7785 59814 10856 59866
rect 1104 59792 10856 59814
rect 753 59755 811 59761
rect 753 59721 765 59755
rect 799 59752 811 59755
rect 1670 59752 1676 59764
rect 799 59724 1676 59752
rect 799 59721 811 59724
rect 753 59715 811 59721
rect 1670 59712 1676 59724
rect 1728 59712 1734 59764
rect 2866 59712 2872 59764
rect 2924 59752 2930 59764
rect 3142 59752 3148 59764
rect 2924 59724 3148 59752
rect 2924 59712 2930 59724
rect 3142 59712 3148 59724
rect 3200 59712 3206 59764
rect 934 59644 940 59696
rect 992 59684 998 59696
rect 992 59656 2176 59684
rect 992 59644 998 59656
rect 1486 59576 1492 59628
rect 1544 59616 1550 59628
rect 2148 59625 2176 59656
rect 1673 59619 1731 59625
rect 1673 59616 1685 59619
rect 1544 59588 1685 59616
rect 1544 59576 1550 59588
rect 1673 59585 1685 59588
rect 1719 59585 1731 59619
rect 1673 59579 1731 59585
rect 2133 59619 2191 59625
rect 2133 59585 2145 59619
rect 2179 59585 2191 59619
rect 2133 59579 2191 59585
rect 1394 59508 1400 59560
rect 1452 59508 1458 59560
rect 1412 59480 1440 59508
rect 2317 59483 2375 59489
rect 2317 59480 2329 59483
rect 1412 59452 2329 59480
rect 2317 59449 2329 59452
rect 2363 59449 2375 59483
rect 2317 59443 2375 59449
rect 842 59372 848 59424
rect 900 59412 906 59424
rect 1489 59415 1547 59421
rect 1489 59412 1501 59415
rect 900 59384 1501 59412
rect 900 59372 906 59384
rect 1489 59381 1501 59384
rect 1535 59381 1547 59415
rect 1489 59375 1547 59381
rect 1104 59322 10856 59344
rect 1104 59270 2582 59322
rect 2634 59270 2646 59322
rect 2698 59270 2710 59322
rect 2762 59270 2774 59322
rect 2826 59270 2838 59322
rect 2890 59270 5845 59322
rect 5897 59270 5909 59322
rect 5961 59270 5973 59322
rect 6025 59270 6037 59322
rect 6089 59270 6101 59322
rect 6153 59270 9109 59322
rect 9161 59270 9173 59322
rect 9225 59270 9237 59322
rect 9289 59270 9301 59322
rect 9353 59270 9365 59322
rect 9417 59270 10856 59322
rect 1104 59248 10856 59270
rect 9858 59168 9864 59220
rect 9916 59208 9922 59220
rect 9953 59211 10011 59217
rect 9953 59208 9965 59211
rect 9916 59180 9965 59208
rect 9916 59168 9922 59180
rect 9953 59177 9965 59180
rect 9999 59177 10011 59211
rect 9953 59171 10011 59177
rect 845 59075 903 59081
rect 845 59041 857 59075
rect 891 59072 903 59075
rect 891 59044 1808 59072
rect 891 59041 903 59044
rect 845 59035 903 59041
rect 750 58964 756 59016
rect 808 59004 814 59016
rect 1673 59007 1731 59013
rect 1673 59004 1685 59007
rect 808 58976 1685 59004
rect 808 58964 814 58976
rect 1673 58973 1685 58976
rect 1719 58973 1731 59007
rect 1780 59004 1808 59044
rect 1854 59032 1860 59084
rect 1912 59072 1918 59084
rect 2409 59075 2467 59081
rect 2409 59072 2421 59075
rect 1912 59044 2421 59072
rect 1912 59032 1918 59044
rect 2409 59041 2421 59044
rect 2455 59041 2467 59075
rect 2409 59035 2467 59041
rect 2133 59007 2191 59013
rect 2133 59004 2145 59007
rect 1780 58976 2145 59004
rect 1673 58967 1731 58973
rect 2133 58973 2145 58976
rect 2179 58973 2191 59007
rect 10134 59004 10140 59016
rect 10095 58976 10140 59004
rect 2133 58967 2191 58973
rect 10134 58964 10140 58976
rect 10192 58964 10198 59016
rect 1486 58868 1492 58880
rect 1447 58840 1492 58868
rect 1486 58828 1492 58840
rect 1544 58828 1550 58880
rect 1104 58778 10856 58800
rect 1104 58726 4213 58778
rect 4265 58726 4277 58778
rect 4329 58726 4341 58778
rect 4393 58726 4405 58778
rect 4457 58726 4469 58778
rect 4521 58726 7477 58778
rect 7529 58726 7541 58778
rect 7593 58726 7605 58778
rect 7657 58726 7669 58778
rect 7721 58726 7733 58778
rect 7785 58726 10856 58778
rect 1104 58704 10856 58726
rect 842 58488 848 58540
rect 900 58528 906 58540
rect 1673 58531 1731 58537
rect 1673 58528 1685 58531
rect 900 58500 1685 58528
rect 900 58488 906 58500
rect 1673 58497 1685 58500
rect 1719 58497 1731 58531
rect 10134 58528 10140 58540
rect 10095 58500 10140 58528
rect 1673 58491 1731 58497
rect 10134 58488 10140 58500
rect 10192 58488 10198 58540
rect 1394 58284 1400 58336
rect 1452 58324 1458 58336
rect 1489 58327 1547 58333
rect 1489 58324 1501 58327
rect 1452 58296 1501 58324
rect 1452 58284 1458 58296
rect 1489 58293 1501 58296
rect 1535 58293 1547 58327
rect 9950 58324 9956 58336
rect 9911 58296 9956 58324
rect 1489 58287 1547 58293
rect 9950 58284 9956 58296
rect 10008 58284 10014 58336
rect 1104 58234 10856 58256
rect 1104 58182 2582 58234
rect 2634 58182 2646 58234
rect 2698 58182 2710 58234
rect 2762 58182 2774 58234
rect 2826 58182 2838 58234
rect 2890 58182 5845 58234
rect 5897 58182 5909 58234
rect 5961 58182 5973 58234
rect 6025 58182 6037 58234
rect 6089 58182 6101 58234
rect 6153 58182 9109 58234
rect 9161 58182 9173 58234
rect 9225 58182 9237 58234
rect 9289 58182 9301 58234
rect 9353 58182 9365 58234
rect 9417 58182 10856 58234
rect 1104 58160 10856 58182
rect 1854 58012 1860 58064
rect 1912 58012 1918 58064
rect 1949 58055 2007 58061
rect 1949 58021 1961 58055
rect 1995 58052 2007 58055
rect 2866 58052 2872 58064
rect 1995 58024 2872 58052
rect 1995 58021 2007 58024
rect 1949 58015 2007 58021
rect 2866 58012 2872 58024
rect 2924 58012 2930 58064
rect 1486 57984 1492 57996
rect 1399 57956 1492 57984
rect 1412 57925 1440 57956
rect 1486 57944 1492 57956
rect 1544 57984 1550 57996
rect 1872 57984 1900 58012
rect 1544 57956 1900 57984
rect 1544 57944 1550 57956
rect 1397 57919 1455 57925
rect 1397 57885 1409 57919
rect 1443 57885 1455 57919
rect 1397 57879 1455 57885
rect 1817 57919 1875 57925
rect 1817 57885 1829 57919
rect 1863 57916 1875 57919
rect 1946 57916 1952 57928
rect 1863 57888 1952 57916
rect 1863 57885 1875 57888
rect 1817 57879 1875 57885
rect 1946 57876 1952 57888
rect 2004 57876 2010 57928
rect 2777 57919 2835 57925
rect 2777 57885 2789 57919
rect 2823 57916 2835 57919
rect 4706 57916 4712 57928
rect 2823 57888 4712 57916
rect 2823 57885 2835 57888
rect 2777 57879 2835 57885
rect 4706 57876 4712 57888
rect 4764 57876 4770 57928
rect 10134 57916 10140 57928
rect 10095 57888 10140 57916
rect 10134 57876 10140 57888
rect 10192 57876 10198 57928
rect 1581 57851 1639 57857
rect 1581 57817 1593 57851
rect 1627 57817 1639 57851
rect 1581 57811 1639 57817
rect 1673 57851 1731 57857
rect 1673 57817 1685 57851
rect 1719 57848 1731 57851
rect 1719 57820 9996 57848
rect 1719 57817 1731 57820
rect 1673 57811 1731 57817
rect 1118 57740 1124 57792
rect 1176 57780 1182 57792
rect 1302 57780 1308 57792
rect 1176 57752 1308 57780
rect 1176 57740 1182 57752
rect 1302 57740 1308 57752
rect 1360 57740 1366 57792
rect 1596 57780 1624 57811
rect 2130 57780 2136 57792
rect 1596 57752 2136 57780
rect 2130 57740 2136 57752
rect 2188 57740 2194 57792
rect 2593 57783 2651 57789
rect 2593 57749 2605 57783
rect 2639 57780 2651 57783
rect 2774 57780 2780 57792
rect 2639 57752 2780 57780
rect 2639 57749 2651 57752
rect 2593 57743 2651 57749
rect 2774 57740 2780 57752
rect 2832 57740 2838 57792
rect 9968 57789 9996 57820
rect 9953 57783 10011 57789
rect 9953 57749 9965 57783
rect 9999 57749 10011 57783
rect 9953 57743 10011 57749
rect 1104 57690 10856 57712
rect 1104 57638 4213 57690
rect 4265 57638 4277 57690
rect 4329 57638 4341 57690
rect 4393 57638 4405 57690
rect 4457 57638 4469 57690
rect 4521 57638 7477 57690
rect 7529 57638 7541 57690
rect 7593 57638 7605 57690
rect 7657 57638 7669 57690
rect 7721 57638 7733 57690
rect 7785 57638 10856 57690
rect 1104 57616 10856 57638
rect 1670 57536 1676 57588
rect 1728 57576 1734 57588
rect 2130 57576 2136 57588
rect 1728 57548 2136 57576
rect 1728 57536 1734 57548
rect 2130 57536 2136 57548
rect 2188 57536 2194 57588
rect 2406 57536 2412 57588
rect 2464 57536 2470 57588
rect 2501 57579 2559 57585
rect 2501 57545 2513 57579
rect 2547 57576 2559 57579
rect 7190 57576 7196 57588
rect 2547 57548 7196 57576
rect 2547 57545 2559 57548
rect 2501 57539 2559 57545
rect 7190 57536 7196 57548
rect 7248 57536 7254 57588
rect 1118 57468 1124 57520
rect 1176 57508 1182 57520
rect 1581 57511 1639 57517
rect 1581 57508 1593 57511
rect 1176 57480 1593 57508
rect 1176 57468 1182 57480
rect 1581 57477 1593 57480
rect 1627 57477 1639 57511
rect 2424 57508 2452 57536
rect 2869 57511 2927 57517
rect 2869 57508 2881 57511
rect 2424 57480 2881 57508
rect 1581 57471 1639 57477
rect 2869 57477 2881 57480
rect 2915 57477 2927 57511
rect 11241 57511 11299 57517
rect 11241 57508 11253 57511
rect 2869 57471 2927 57477
rect 2976 57480 11253 57508
rect 1397 57443 1455 57449
rect 1397 57409 1409 57443
rect 1443 57440 1455 57443
rect 1486 57440 1492 57452
rect 1443 57412 1492 57440
rect 1443 57409 1455 57412
rect 1397 57403 1455 57409
rect 1486 57400 1492 57412
rect 1544 57400 1550 57452
rect 1673 57443 1731 57449
rect 1673 57409 1685 57443
rect 1719 57409 1731 57443
rect 1673 57403 1731 57409
rect 1817 57443 1875 57449
rect 1817 57409 1829 57443
rect 1863 57440 1875 57443
rect 1946 57440 1952 57452
rect 1863 57412 1952 57440
rect 1863 57409 1875 57412
rect 1817 57403 1875 57409
rect 1688 57372 1716 57403
rect 1946 57400 1952 57412
rect 2004 57400 2010 57452
rect 2314 57400 2320 57452
rect 2372 57440 2378 57452
rect 2685 57443 2743 57449
rect 2685 57440 2697 57443
rect 2372 57412 2697 57440
rect 2372 57400 2378 57412
rect 2685 57409 2697 57412
rect 2731 57409 2743 57443
rect 2685 57403 2743 57409
rect 2777 57443 2835 57449
rect 2777 57409 2789 57443
rect 2823 57440 2835 57443
rect 2976 57440 3004 57480
rect 11241 57477 11253 57480
rect 11287 57477 11299 57511
rect 11241 57471 11299 57477
rect 2823 57412 3004 57440
rect 3053 57443 3111 57449
rect 2823 57409 2835 57412
rect 2777 57403 2835 57409
rect 3053 57409 3065 57443
rect 3099 57440 3111 57443
rect 3326 57440 3332 57452
rect 3099 57412 3332 57440
rect 3099 57409 3111 57412
rect 3053 57403 3111 57409
rect 3326 57400 3332 57412
rect 3384 57400 3390 57452
rect 9950 57372 9956 57384
rect 1688 57344 9956 57372
rect 9950 57332 9956 57344
rect 10008 57332 10014 57384
rect 1949 57307 2007 57313
rect 1949 57273 1961 57307
rect 1995 57304 2007 57307
rect 3694 57304 3700 57316
rect 1995 57276 3700 57304
rect 1995 57273 2007 57276
rect 1949 57267 2007 57273
rect 3694 57264 3700 57276
rect 3752 57264 3758 57316
rect 1670 57196 1676 57248
rect 1728 57236 1734 57248
rect 5442 57236 5448 57248
rect 1728 57208 5448 57236
rect 1728 57196 1734 57208
rect 5442 57196 5448 57208
rect 5500 57196 5506 57248
rect 1104 57146 10856 57168
rect 1104 57094 2582 57146
rect 2634 57094 2646 57146
rect 2698 57094 2710 57146
rect 2762 57094 2774 57146
rect 2826 57094 2838 57146
rect 2890 57094 5845 57146
rect 5897 57094 5909 57146
rect 5961 57094 5973 57146
rect 6025 57094 6037 57146
rect 6089 57094 6101 57146
rect 6153 57094 9109 57146
rect 9161 57094 9173 57146
rect 9225 57094 9237 57146
rect 9289 57094 9301 57146
rect 9353 57094 9365 57146
rect 9417 57094 10856 57146
rect 1104 57072 10856 57094
rect 2314 56924 2320 56976
rect 2372 56964 2378 56976
rect 2372 56936 2728 56964
rect 2372 56924 2378 56936
rect 2590 56856 2596 56908
rect 2648 56856 2654 56908
rect 1670 56828 1676 56840
rect 1631 56800 1676 56828
rect 1670 56788 1676 56800
rect 1728 56788 1734 56840
rect 2317 56831 2375 56837
rect 2317 56797 2329 56831
rect 2363 56828 2375 56831
rect 2608 56828 2636 56856
rect 2700 56837 2728 56936
rect 2774 56924 2780 56976
rect 2832 56964 2838 56976
rect 3326 56964 3332 56976
rect 2832 56936 3332 56964
rect 2832 56924 2838 56936
rect 3326 56924 3332 56936
rect 3384 56924 3390 56976
rect 9861 56899 9919 56905
rect 9861 56865 9873 56899
rect 9907 56896 9919 56899
rect 11701 56899 11759 56905
rect 11701 56896 11713 56899
rect 9907 56868 11713 56896
rect 9907 56865 9919 56868
rect 9861 56859 9919 56865
rect 11701 56865 11713 56868
rect 11747 56865 11759 56899
rect 11701 56859 11759 56865
rect 2363 56800 2636 56828
rect 2685 56831 2743 56837
rect 2363 56797 2375 56800
rect 2317 56791 2375 56797
rect 2685 56797 2697 56831
rect 2731 56797 2743 56831
rect 10134 56828 10140 56840
rect 10095 56800 10140 56828
rect 2685 56791 2743 56797
rect 10134 56788 10140 56800
rect 10192 56788 10198 56840
rect 2498 56760 2504 56772
rect 2459 56732 2504 56760
rect 2498 56720 2504 56732
rect 2556 56720 2562 56772
rect 2593 56763 2651 56769
rect 2593 56729 2605 56763
rect 2639 56760 2651 56763
rect 11425 56763 11483 56769
rect 11425 56760 11437 56763
rect 2639 56732 11437 56760
rect 2639 56729 2651 56732
rect 2593 56723 2651 56729
rect 11425 56729 11437 56732
rect 11471 56729 11483 56763
rect 11425 56723 11483 56729
rect 1486 56692 1492 56704
rect 1447 56664 1492 56692
rect 1486 56652 1492 56664
rect 1544 56652 1550 56704
rect 2869 56695 2927 56701
rect 2869 56661 2881 56695
rect 2915 56692 2927 56695
rect 8754 56692 8760 56704
rect 2915 56664 8760 56692
rect 2915 56661 2927 56664
rect 2869 56655 2927 56661
rect 8754 56652 8760 56664
rect 8812 56652 8818 56704
rect 1104 56602 10856 56624
rect 1104 56550 4213 56602
rect 4265 56550 4277 56602
rect 4329 56550 4341 56602
rect 4393 56550 4405 56602
rect 4457 56550 4469 56602
rect 4521 56550 7477 56602
rect 7529 56550 7541 56602
rect 7593 56550 7605 56602
rect 7657 56550 7669 56602
rect 7721 56550 7733 56602
rect 7785 56550 10856 56602
rect 1104 56528 10856 56550
rect 1394 56448 1400 56500
rect 1452 56488 1458 56500
rect 1489 56491 1547 56497
rect 1489 56488 1501 56491
rect 1452 56460 1501 56488
rect 1452 56448 1458 56460
rect 1489 56457 1501 56460
rect 1535 56457 1547 56491
rect 1489 56451 1547 56457
rect 1670 56448 1676 56500
rect 1728 56488 1734 56500
rect 3602 56488 3608 56500
rect 1728 56460 3608 56488
rect 1728 56448 1734 56460
rect 3602 56448 3608 56460
rect 3660 56448 3666 56500
rect 1854 56380 1860 56432
rect 1912 56420 1918 56432
rect 2314 56420 2320 56432
rect 1912 56392 2320 56420
rect 1912 56380 1918 56392
rect 2314 56380 2320 56392
rect 2372 56380 2378 56432
rect 2409 56423 2467 56429
rect 2409 56389 2421 56423
rect 2455 56420 2467 56423
rect 2774 56420 2780 56432
rect 2455 56392 2780 56420
rect 2455 56389 2467 56392
rect 2409 56383 2467 56389
rect 2774 56380 2780 56392
rect 2832 56380 2838 56432
rect 1673 56355 1731 56361
rect 1673 56321 1685 56355
rect 1719 56352 1731 56355
rect 2961 56355 3019 56361
rect 1719 56324 2774 56352
rect 1719 56321 1731 56324
rect 1673 56315 1731 56321
rect 2746 56284 2774 56324
rect 2961 56321 2973 56355
rect 3007 56352 3019 56355
rect 8846 56352 8852 56364
rect 3007 56324 8852 56352
rect 3007 56321 3019 56324
rect 2961 56315 3019 56321
rect 8846 56312 8852 56324
rect 8904 56312 8910 56364
rect 10134 56352 10140 56364
rect 10095 56324 10140 56352
rect 10134 56312 10140 56324
rect 10192 56312 10198 56364
rect 3234 56284 3240 56296
rect 2746 56256 3240 56284
rect 3234 56244 3240 56256
rect 3292 56244 3298 56296
rect 3602 56244 3608 56296
rect 3660 56284 3666 56296
rect 3970 56284 3976 56296
rect 3660 56256 3976 56284
rect 3660 56244 3666 56256
rect 3970 56244 3976 56256
rect 4028 56244 4034 56296
rect 1854 56176 1860 56228
rect 1912 56216 1918 56228
rect 2225 56219 2283 56225
rect 2225 56216 2237 56219
rect 1912 56188 2237 56216
rect 1912 56176 1918 56188
rect 2225 56185 2237 56188
rect 2271 56185 2283 56219
rect 2225 56179 2283 56185
rect 2866 56176 2872 56228
rect 2924 56216 2930 56228
rect 3050 56216 3056 56228
rect 2924 56188 3056 56216
rect 2924 56176 2930 56188
rect 3050 56176 3056 56188
rect 3108 56176 3114 56228
rect 3142 56148 3148 56160
rect 3103 56120 3148 56148
rect 3142 56108 3148 56120
rect 3200 56108 3206 56160
rect 9950 56148 9956 56160
rect 9911 56120 9956 56148
rect 9950 56108 9956 56120
rect 10008 56108 10014 56160
rect 1104 56058 10856 56080
rect 1104 56006 2582 56058
rect 2634 56006 2646 56058
rect 2698 56006 2710 56058
rect 2762 56006 2774 56058
rect 2826 56006 2838 56058
rect 2890 56006 5845 56058
rect 5897 56006 5909 56058
rect 5961 56006 5973 56058
rect 6025 56006 6037 56058
rect 6089 56006 6101 56058
rect 6153 56006 9109 56058
rect 9161 56006 9173 56058
rect 9225 56006 9237 56058
rect 9289 56006 9301 56058
rect 9353 56006 9365 56058
rect 9417 56006 10856 56058
rect 1104 55984 10856 56006
rect 937 55947 995 55953
rect 937 55913 949 55947
rect 983 55944 995 55947
rect 2406 55944 2412 55956
rect 983 55916 2412 55944
rect 983 55913 995 55916
rect 937 55907 995 55913
rect 2406 55904 2412 55916
rect 2464 55904 2470 55956
rect 3237 55879 3295 55885
rect 3237 55845 3249 55879
rect 3283 55876 3295 55879
rect 3326 55876 3332 55888
rect 3283 55848 3332 55876
rect 3283 55845 3295 55848
rect 3237 55839 3295 55845
rect 3326 55836 3332 55848
rect 3384 55836 3390 55888
rect 7926 55808 7932 55820
rect 1688 55780 7932 55808
rect 1688 55749 1716 55780
rect 7926 55768 7932 55780
rect 7984 55768 7990 55820
rect 1673 55743 1731 55749
rect 1673 55709 1685 55743
rect 1719 55709 1731 55743
rect 1673 55703 1731 55709
rect 2225 55743 2283 55749
rect 2225 55709 2237 55743
rect 2271 55740 2283 55743
rect 3789 55743 3847 55749
rect 2271 55712 3096 55740
rect 2271 55709 2283 55712
rect 2225 55703 2283 55709
rect 3068 55681 3096 55712
rect 3789 55709 3801 55743
rect 3835 55740 3847 55743
rect 8662 55740 8668 55752
rect 3835 55712 8668 55740
rect 3835 55709 3847 55712
rect 3789 55703 3847 55709
rect 8662 55700 8668 55712
rect 8720 55700 8726 55752
rect 10965 55743 11023 55749
rect 10965 55709 10977 55743
rect 11011 55740 11023 55743
rect 11517 55743 11575 55749
rect 11517 55740 11529 55743
rect 11011 55712 11529 55740
rect 11011 55709 11023 55712
rect 10965 55703 11023 55709
rect 11517 55709 11529 55712
rect 11563 55709 11575 55743
rect 11517 55703 11575 55709
rect 845 55675 903 55681
rect 845 55641 857 55675
rect 891 55672 903 55675
rect 3053 55675 3111 55681
rect 891 55644 2452 55672
rect 891 55641 903 55644
rect 845 55635 903 55641
rect 1486 55604 1492 55616
rect 1447 55576 1492 55604
rect 1486 55564 1492 55576
rect 1544 55564 1550 55616
rect 2424 55613 2452 55644
rect 3053 55641 3065 55675
rect 3099 55672 3111 55675
rect 3142 55672 3148 55684
rect 3099 55644 3148 55672
rect 3099 55641 3111 55644
rect 3053 55635 3111 55641
rect 3142 55632 3148 55644
rect 3200 55632 3206 55684
rect 11885 55675 11943 55681
rect 11885 55672 11897 55675
rect 3252 55644 11897 55672
rect 2409 55607 2467 55613
rect 2409 55573 2421 55607
rect 2455 55604 2467 55607
rect 2498 55604 2504 55616
rect 2455 55576 2504 55604
rect 2455 55573 2467 55576
rect 2409 55567 2467 55573
rect 2498 55564 2504 55576
rect 2556 55564 2562 55616
rect 2774 55564 2780 55616
rect 2832 55604 2838 55616
rect 3252 55604 3280 55644
rect 11885 55641 11897 55644
rect 11931 55641 11943 55675
rect 11885 55635 11943 55641
rect 3970 55604 3976 55616
rect 2832 55576 3280 55604
rect 3931 55576 3976 55604
rect 2832 55564 2838 55576
rect 3970 55564 3976 55576
rect 4028 55564 4034 55616
rect 1104 55514 10856 55536
rect 1104 55462 4213 55514
rect 4265 55462 4277 55514
rect 4329 55462 4341 55514
rect 4393 55462 4405 55514
rect 4457 55462 4469 55514
rect 4521 55462 7477 55514
rect 7529 55462 7541 55514
rect 7593 55462 7605 55514
rect 7657 55462 7669 55514
rect 7721 55462 7733 55514
rect 7785 55462 10856 55514
rect 1104 55440 10856 55462
rect 9950 55400 9956 55412
rect 1688 55372 9956 55400
rect 1688 55341 1716 55372
rect 9950 55360 9956 55372
rect 10008 55360 10014 55412
rect 1673 55335 1731 55341
rect 1673 55301 1685 55335
rect 1719 55301 1731 55335
rect 1673 55295 1731 55301
rect 1966 55335 2024 55341
rect 1966 55301 1978 55335
rect 2012 55332 2024 55335
rect 2774 55332 2780 55344
rect 2012 55304 2780 55332
rect 2012 55301 2024 55304
rect 1966 55295 2024 55301
rect 2774 55292 2780 55304
rect 2832 55292 2838 55344
rect 3234 55292 3240 55344
rect 3292 55332 3298 55344
rect 3970 55332 3976 55344
rect 3292 55304 3976 55332
rect 3292 55292 3298 55304
rect 3970 55292 3976 55304
rect 4028 55292 4034 55344
rect 1854 55273 1860 55276
rect 1397 55267 1455 55273
rect 1397 55233 1409 55267
rect 1443 55233 1455 55267
rect 1397 55227 1455 55233
rect 1581 55267 1639 55273
rect 1581 55233 1593 55267
rect 1627 55264 1639 55267
rect 1817 55267 1860 55273
rect 1627 55236 1716 55264
rect 1627 55233 1639 55236
rect 1581 55227 1639 55233
rect 1412 55060 1440 55227
rect 1688 55208 1716 55236
rect 1817 55233 1829 55267
rect 1817 55227 1860 55233
rect 1854 55224 1860 55227
rect 1912 55224 1918 55276
rect 2501 55267 2559 55273
rect 2501 55233 2513 55267
rect 2547 55264 2559 55267
rect 8386 55264 8392 55276
rect 2547 55236 8392 55264
rect 2547 55233 2559 55236
rect 2501 55227 2559 55233
rect 8386 55224 8392 55236
rect 8444 55224 8450 55276
rect 10134 55264 10140 55276
rect 10095 55236 10140 55264
rect 10134 55224 10140 55236
rect 10192 55224 10198 55276
rect 1670 55156 1676 55208
rect 1728 55156 1734 55208
rect 2685 55131 2743 55137
rect 2685 55097 2697 55131
rect 2731 55128 2743 55131
rect 2774 55128 2780 55140
rect 2731 55100 2780 55128
rect 2731 55097 2743 55100
rect 2685 55091 2743 55097
rect 2774 55088 2780 55100
rect 2832 55088 2838 55140
rect 1670 55060 1676 55072
rect 1412 55032 1676 55060
rect 1670 55020 1676 55032
rect 1728 55020 1734 55072
rect 9950 55060 9956 55072
rect 9911 55032 9956 55060
rect 9950 55020 9956 55032
rect 10008 55020 10014 55072
rect 1104 54970 10856 54992
rect 1104 54918 2582 54970
rect 2634 54918 2646 54970
rect 2698 54918 2710 54970
rect 2762 54918 2774 54970
rect 2826 54918 2838 54970
rect 2890 54918 5845 54970
rect 5897 54918 5909 54970
rect 5961 54918 5973 54970
rect 6025 54918 6037 54970
rect 6089 54918 6101 54970
rect 6153 54918 9109 54970
rect 9161 54918 9173 54970
rect 9225 54918 9237 54970
rect 9289 54918 9301 54970
rect 9353 54918 9365 54970
rect 9417 54918 10856 54970
rect 1104 54896 10856 54918
rect 1673 54655 1731 54661
rect 1673 54621 1685 54655
rect 1719 54621 1731 54655
rect 1673 54615 1731 54621
rect 2409 54655 2467 54661
rect 2409 54621 2421 54655
rect 2455 54652 2467 54655
rect 6822 54652 6828 54664
rect 2455 54624 6828 54652
rect 2455 54621 2467 54624
rect 2409 54615 2467 54621
rect 1688 54584 1716 54615
rect 6822 54612 6828 54624
rect 6880 54612 6886 54664
rect 10134 54652 10140 54664
rect 10095 54624 10140 54652
rect 10134 54612 10140 54624
rect 10192 54612 10198 54664
rect 7282 54584 7288 54596
rect 1688 54556 7288 54584
rect 7282 54544 7288 54556
rect 7340 54544 7346 54596
rect 1486 54516 1492 54528
rect 1447 54488 1492 54516
rect 1486 54476 1492 54488
rect 1544 54476 1550 54528
rect 2222 54516 2228 54528
rect 2183 54488 2228 54516
rect 2222 54476 2228 54488
rect 2280 54476 2286 54528
rect 9953 54519 10011 54525
rect 9953 54485 9965 54519
rect 9999 54516 10011 54519
rect 10965 54519 11023 54525
rect 10965 54516 10977 54519
rect 9999 54488 10977 54516
rect 9999 54485 10011 54488
rect 9953 54479 10011 54485
rect 10965 54485 10977 54488
rect 11011 54485 11023 54519
rect 10965 54479 11023 54485
rect 1104 54426 10856 54448
rect 1104 54374 4213 54426
rect 4265 54374 4277 54426
rect 4329 54374 4341 54426
rect 4393 54374 4405 54426
rect 4457 54374 4469 54426
rect 4521 54374 7477 54426
rect 7529 54374 7541 54426
rect 7593 54374 7605 54426
rect 7657 54374 7669 54426
rect 7721 54374 7733 54426
rect 7785 54374 10856 54426
rect 1104 54352 10856 54374
rect 2961 54315 3019 54321
rect 2961 54281 2973 54315
rect 3007 54312 3019 54315
rect 3050 54312 3056 54324
rect 3007 54284 3056 54312
rect 3007 54281 3019 54284
rect 2961 54275 3019 54281
rect 3050 54272 3056 54284
rect 3108 54272 3114 54324
rect 1581 54179 1639 54185
rect 1581 54145 1593 54179
rect 1627 54176 1639 54179
rect 2498 54176 2504 54188
rect 1627 54148 2504 54176
rect 1627 54145 1639 54148
rect 1581 54139 1639 54145
rect 2498 54136 2504 54148
rect 2556 54136 2562 54188
rect 2869 54179 2927 54185
rect 2869 54145 2881 54179
rect 2915 54176 2927 54179
rect 2958 54176 2964 54188
rect 2915 54148 2964 54176
rect 2915 54145 2927 54148
rect 2869 54139 2927 54145
rect 2958 54136 2964 54148
rect 3016 54136 3022 54188
rect 3053 54179 3111 54185
rect 3053 54145 3065 54179
rect 3099 54176 3111 54179
rect 3326 54176 3332 54188
rect 3099 54148 3332 54176
rect 3099 54145 3111 54148
rect 3053 54139 3111 54145
rect 3326 54136 3332 54148
rect 3384 54136 3390 54188
rect 5718 54136 5724 54188
rect 5776 54176 5782 54188
rect 6270 54176 6276 54188
rect 5776 54148 6276 54176
rect 5776 54136 5782 54148
rect 6270 54136 6276 54148
rect 6328 54136 6334 54188
rect 9766 54136 9772 54188
rect 9824 54176 9830 54188
rect 9861 54179 9919 54185
rect 9861 54176 9873 54179
rect 9824 54148 9873 54176
rect 9824 54136 9830 54148
rect 9861 54145 9873 54148
rect 9907 54145 9919 54179
rect 9861 54139 9919 54145
rect 11241 54179 11299 54185
rect 11241 54145 11253 54179
rect 11287 54176 11299 54179
rect 11609 54179 11667 54185
rect 11609 54176 11621 54179
rect 11287 54148 11621 54176
rect 11287 54145 11299 54148
rect 11241 54139 11299 54145
rect 11609 54145 11621 54148
rect 11655 54145 11667 54179
rect 11609 54139 11667 54145
rect 1670 54068 1676 54120
rect 1728 54108 1734 54120
rect 1857 54111 1915 54117
rect 1857 54108 1869 54111
rect 1728 54080 1869 54108
rect 1728 54068 1734 54080
rect 1857 54077 1869 54080
rect 1903 54077 1915 54111
rect 1857 54071 1915 54077
rect 10042 53972 10048 53984
rect 10003 53944 10048 53972
rect 10042 53932 10048 53944
rect 10100 53932 10106 53984
rect 11517 53975 11575 53981
rect 11517 53941 11529 53975
rect 11563 53972 11575 53975
rect 11701 53975 11759 53981
rect 11701 53972 11713 53975
rect 11563 53944 11713 53972
rect 11563 53941 11575 53944
rect 11517 53935 11575 53941
rect 11701 53941 11713 53944
rect 11747 53941 11759 53975
rect 11701 53935 11759 53941
rect 1104 53882 10856 53904
rect 1104 53830 2582 53882
rect 2634 53830 2646 53882
rect 2698 53830 2710 53882
rect 2762 53830 2774 53882
rect 2826 53830 2838 53882
rect 2890 53830 5845 53882
rect 5897 53830 5909 53882
rect 5961 53830 5973 53882
rect 6025 53830 6037 53882
rect 6089 53830 6101 53882
rect 6153 53830 9109 53882
rect 9161 53830 9173 53882
rect 9225 53830 9237 53882
rect 9289 53830 9301 53882
rect 9353 53830 9365 53882
rect 9417 53830 10856 53882
rect 1104 53808 10856 53830
rect 1762 53660 1768 53712
rect 1820 53660 1826 53712
rect 1949 53703 2007 53709
rect 1949 53669 1961 53703
rect 1995 53700 2007 53703
rect 11701 53703 11759 53709
rect 11701 53700 11713 53703
rect 1995 53672 11713 53700
rect 1995 53669 2007 53672
rect 1949 53663 2007 53669
rect 11701 53669 11713 53672
rect 11747 53669 11759 53703
rect 11701 53663 11759 53669
rect 1780 53632 1808 53660
rect 1596 53604 1808 53632
rect 1397 53567 1455 53573
rect 1397 53533 1409 53567
rect 1443 53564 1455 53567
rect 1486 53564 1492 53576
rect 1443 53536 1492 53564
rect 1443 53533 1455 53536
rect 1397 53527 1455 53533
rect 1486 53524 1492 53536
rect 1544 53524 1550 53576
rect 1596 53573 1624 53604
rect 1854 53573 1860 53576
rect 1581 53567 1639 53573
rect 1581 53533 1593 53567
rect 1627 53533 1639 53567
rect 1581 53527 1639 53533
rect 1817 53567 1860 53573
rect 1817 53533 1829 53567
rect 1817 53527 1860 53533
rect 1854 53524 1860 53527
rect 1912 53524 1918 53576
rect 2501 53567 2559 53573
rect 2501 53533 2513 53567
rect 2547 53564 2559 53567
rect 8018 53564 8024 53576
rect 2547 53536 8024 53564
rect 2547 53533 2559 53536
rect 2501 53527 2559 53533
rect 8018 53524 8024 53536
rect 8076 53524 8082 53576
rect 1673 53499 1731 53505
rect 1673 53465 1685 53499
rect 1719 53496 1731 53499
rect 9950 53496 9956 53508
rect 1719 53468 9956 53496
rect 1719 53465 1731 53468
rect 1673 53459 1731 53465
rect 9950 53456 9956 53468
rect 10008 53456 10014 53508
rect 1762 53388 1768 53440
rect 1820 53428 1826 53440
rect 2130 53428 2136 53440
rect 1820 53400 2136 53428
rect 1820 53388 1826 53400
rect 2130 53388 2136 53400
rect 2188 53388 2194 53440
rect 2685 53431 2743 53437
rect 2685 53397 2697 53431
rect 2731 53428 2743 53431
rect 2774 53428 2780 53440
rect 2731 53400 2780 53428
rect 2731 53397 2743 53400
rect 2685 53391 2743 53397
rect 2774 53388 2780 53400
rect 2832 53388 2838 53440
rect 1104 53338 10856 53360
rect 1104 53286 4213 53338
rect 4265 53286 4277 53338
rect 4329 53286 4341 53338
rect 4393 53286 4405 53338
rect 4457 53286 4469 53338
rect 4521 53286 7477 53338
rect 7529 53286 7541 53338
rect 7593 53286 7605 53338
rect 7657 53286 7669 53338
rect 7721 53286 7733 53338
rect 7785 53286 10856 53338
rect 1104 53264 10856 53286
rect 1486 53184 1492 53236
rect 1544 53224 1550 53236
rect 1670 53224 1676 53236
rect 1544 53196 1676 53224
rect 1544 53184 1550 53196
rect 1670 53184 1676 53196
rect 1728 53224 1734 53236
rect 2498 53224 2504 53236
rect 1728 53196 2504 53224
rect 1728 53184 1734 53196
rect 2498 53184 2504 53196
rect 2556 53184 2562 53236
rect 6638 53156 6644 53168
rect 2746 53128 6644 53156
rect 1673 53091 1731 53097
rect 1673 53057 1685 53091
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 2409 53091 2467 53097
rect 2409 53057 2421 53091
rect 2455 53088 2467 53091
rect 2746 53088 2774 53128
rect 6638 53116 6644 53128
rect 6696 53116 6702 53168
rect 2455 53060 2774 53088
rect 2869 53091 2927 53097
rect 2455 53057 2467 53060
rect 2409 53051 2467 53057
rect 2869 53057 2881 53091
rect 2915 53088 2927 53091
rect 8110 53088 8116 53100
rect 2915 53060 8116 53088
rect 2915 53057 2927 53060
rect 2869 53051 2927 53057
rect 1688 53020 1716 53051
rect 8110 53048 8116 53060
rect 8168 53048 8174 53100
rect 9858 53088 9864 53100
rect 9819 53060 9864 53088
rect 9858 53048 9864 53060
rect 9916 53048 9922 53100
rect 5258 53020 5264 53032
rect 1688 52992 5264 53020
rect 5258 52980 5264 52992
rect 5316 52980 5322 53032
rect 3050 52952 3056 52964
rect 3011 52924 3056 52952
rect 3050 52912 3056 52924
rect 3108 52912 3114 52964
rect 1394 52844 1400 52896
rect 1452 52884 1458 52896
rect 1489 52887 1547 52893
rect 1489 52884 1501 52887
rect 1452 52856 1501 52884
rect 1452 52844 1458 52856
rect 1489 52853 1501 52856
rect 1535 52853 1547 52887
rect 2222 52884 2228 52896
rect 2183 52856 2228 52884
rect 1489 52847 1547 52853
rect 2222 52844 2228 52856
rect 2280 52844 2286 52896
rect 10042 52884 10048 52896
rect 10003 52856 10048 52884
rect 10042 52844 10048 52856
rect 10100 52844 10106 52896
rect 1104 52794 10856 52816
rect 1104 52742 2582 52794
rect 2634 52742 2646 52794
rect 2698 52742 2710 52794
rect 2762 52742 2774 52794
rect 2826 52742 2838 52794
rect 2890 52742 5845 52794
rect 5897 52742 5909 52794
rect 5961 52742 5973 52794
rect 6025 52742 6037 52794
rect 6089 52742 6101 52794
rect 6153 52742 9109 52794
rect 9161 52742 9173 52794
rect 9225 52742 9237 52794
rect 9289 52742 9301 52794
rect 9353 52742 9365 52794
rect 9417 52742 10856 52794
rect 1104 52720 10856 52742
rect 2133 52683 2191 52689
rect 2133 52649 2145 52683
rect 2179 52680 2191 52683
rect 2406 52680 2412 52692
rect 2179 52652 2412 52680
rect 2179 52649 2191 52652
rect 2133 52643 2191 52649
rect 2406 52640 2412 52652
rect 2464 52640 2470 52692
rect 2961 52683 3019 52689
rect 2961 52649 2973 52683
rect 3007 52680 3019 52683
rect 9766 52680 9772 52692
rect 3007 52652 9772 52680
rect 3007 52649 3019 52652
rect 2961 52643 3019 52649
rect 9766 52640 9772 52652
rect 9824 52640 9830 52692
rect 2240 52516 2820 52544
rect 2240 52488 2268 52516
rect 1210 52436 1216 52488
rect 1268 52476 1274 52488
rect 1673 52479 1731 52485
rect 1673 52476 1685 52479
rect 1268 52448 1685 52476
rect 1268 52436 1274 52448
rect 1673 52445 1685 52448
rect 1719 52445 1731 52479
rect 1673 52439 1731 52445
rect 2133 52479 2191 52485
rect 2133 52445 2145 52479
rect 2179 52445 2191 52479
rect 2133 52439 2191 52445
rect 2148 52408 2176 52439
rect 2222 52436 2228 52488
rect 2280 52436 2286 52488
rect 2317 52479 2375 52485
rect 2317 52445 2329 52479
rect 2363 52476 2375 52479
rect 2406 52476 2412 52488
rect 2363 52448 2412 52476
rect 2363 52445 2375 52448
rect 2317 52439 2375 52445
rect 2406 52436 2412 52448
rect 2464 52436 2470 52488
rect 2792 52485 2820 52516
rect 2777 52479 2835 52485
rect 2777 52445 2789 52479
rect 2823 52445 2835 52479
rect 2777 52439 2835 52445
rect 2961 52479 3019 52485
rect 2961 52445 2973 52479
rect 3007 52476 3019 52479
rect 3050 52476 3056 52488
rect 3007 52448 3056 52476
rect 3007 52445 3019 52448
rect 2961 52439 3019 52445
rect 3050 52436 3056 52448
rect 3108 52436 3114 52488
rect 9861 52479 9919 52485
rect 9861 52445 9873 52479
rect 9907 52445 9919 52479
rect 9861 52439 9919 52445
rect 2866 52408 2872 52420
rect 2148 52380 2872 52408
rect 2866 52368 2872 52380
rect 2924 52368 2930 52420
rect 3142 52368 3148 52420
rect 3200 52408 3206 52420
rect 9876 52408 9904 52439
rect 3200 52380 9904 52408
rect 3200 52368 3206 52380
rect 1486 52340 1492 52352
rect 1447 52312 1492 52340
rect 1486 52300 1492 52312
rect 1544 52300 1550 52352
rect 2314 52300 2320 52352
rect 2372 52340 2378 52352
rect 7374 52340 7380 52352
rect 2372 52312 7380 52340
rect 2372 52300 2378 52312
rect 7374 52300 7380 52312
rect 7432 52300 7438 52352
rect 10042 52340 10048 52352
rect 10003 52312 10048 52340
rect 10042 52300 10048 52312
rect 10100 52300 10106 52352
rect 1104 52250 10856 52272
rect 1104 52198 4213 52250
rect 4265 52198 4277 52250
rect 4329 52198 4341 52250
rect 4393 52198 4405 52250
rect 4457 52198 4469 52250
rect 4521 52198 7477 52250
rect 7529 52198 7541 52250
rect 7593 52198 7605 52250
rect 7657 52198 7669 52250
rect 7721 52198 7733 52250
rect 7785 52198 10856 52250
rect 1104 52176 10856 52198
rect 2961 52139 3019 52145
rect 2961 52105 2973 52139
rect 3007 52136 3019 52139
rect 3142 52136 3148 52148
rect 3007 52108 3148 52136
rect 3007 52105 3019 52108
rect 2961 52099 3019 52105
rect 3142 52096 3148 52108
rect 3200 52096 3206 52148
rect 3605 52139 3663 52145
rect 3605 52105 3617 52139
rect 3651 52136 3663 52139
rect 9858 52136 9864 52148
rect 3651 52108 9864 52136
rect 3651 52105 3663 52108
rect 3605 52099 3663 52105
rect 9858 52096 9864 52108
rect 9916 52096 9922 52148
rect 566 52028 572 52080
rect 624 52068 630 52080
rect 624 52040 3740 52068
rect 624 52028 630 52040
rect 1673 52003 1731 52009
rect 1673 51969 1685 52003
rect 1719 52000 1731 52003
rect 2314 52000 2320 52012
rect 1719 51972 2320 52000
rect 1719 51969 1731 51972
rect 1673 51963 1731 51969
rect 2314 51960 2320 51972
rect 2372 51960 2378 52012
rect 2869 52003 2927 52009
rect 2869 51969 2881 52003
rect 2915 52000 2927 52003
rect 2958 52000 2964 52012
rect 2915 51972 2964 52000
rect 2915 51969 2927 51972
rect 2869 51963 2927 51969
rect 2958 51960 2964 51972
rect 3016 51960 3022 52012
rect 3050 51960 3056 52012
rect 3108 52009 3114 52012
rect 3108 52003 3123 52009
rect 3111 52000 3123 52003
rect 3160 52000 3188 52040
rect 3712 52009 3740 52040
rect 3513 52003 3571 52009
rect 3111 51972 3201 52000
rect 3111 51969 3123 51972
rect 3108 51963 3123 51969
rect 3513 51969 3525 52003
rect 3559 51969 3571 52003
rect 3513 51963 3571 51969
rect 3697 52003 3755 52009
rect 3697 51969 3709 52003
rect 3743 51969 3755 52003
rect 3697 51963 3755 51969
rect 3108 51960 3114 51963
rect 937 51935 995 51941
rect 937 51901 949 51935
rect 983 51932 995 51935
rect 3528 51932 3556 51963
rect 983 51904 3556 51932
rect 983 51901 995 51904
rect 937 51895 995 51901
rect 2130 51824 2136 51876
rect 2188 51864 2194 51876
rect 2314 51864 2320 51876
rect 2188 51836 2320 51864
rect 2188 51824 2194 51836
rect 2314 51824 2320 51836
rect 2372 51824 2378 51876
rect 2866 51824 2872 51876
rect 2924 51864 2930 51876
rect 3142 51864 3148 51876
rect 2924 51836 3148 51864
rect 2924 51824 2930 51836
rect 3142 51824 3148 51836
rect 3200 51824 3206 51876
rect 1302 51756 1308 51808
rect 1360 51796 1366 51808
rect 1489 51799 1547 51805
rect 1489 51796 1501 51799
rect 1360 51768 1501 51796
rect 1360 51756 1366 51768
rect 1489 51765 1501 51768
rect 1535 51765 1547 51799
rect 1489 51759 1547 51765
rect 1670 51756 1676 51808
rect 1728 51796 1734 51808
rect 8202 51796 8208 51808
rect 1728 51768 8208 51796
rect 1728 51756 1734 51768
rect 8202 51756 8208 51768
rect 8260 51756 8266 51808
rect 1104 51706 10856 51728
rect 1104 51654 2582 51706
rect 2634 51654 2646 51706
rect 2698 51654 2710 51706
rect 2762 51654 2774 51706
rect 2826 51654 2838 51706
rect 2890 51654 5845 51706
rect 5897 51654 5909 51706
rect 5961 51654 5973 51706
rect 6025 51654 6037 51706
rect 6089 51654 6101 51706
rect 6153 51654 9109 51706
rect 9161 51654 9173 51706
rect 9225 51654 9237 51706
rect 9289 51654 9301 51706
rect 9353 51654 9365 51706
rect 9417 51654 10856 51706
rect 1104 51632 10856 51654
rect 2869 51595 2927 51601
rect 2869 51561 2881 51595
rect 2915 51592 2927 51595
rect 3786 51592 3792 51604
rect 2915 51564 3792 51592
rect 2915 51561 2927 51564
rect 2869 51555 2927 51561
rect 3786 51552 3792 51564
rect 3844 51552 3850 51604
rect 2406 51524 2412 51536
rect 2240 51496 2412 51524
rect 1670 51388 1676 51400
rect 1631 51360 1676 51388
rect 1670 51348 1676 51360
rect 1728 51348 1734 51400
rect 2240 51320 2268 51496
rect 2406 51484 2412 51496
rect 2464 51484 2470 51536
rect 2682 51484 2688 51536
rect 2740 51524 2746 51536
rect 3694 51524 3700 51536
rect 2740 51496 3700 51524
rect 2740 51484 2746 51496
rect 3694 51484 3700 51496
rect 3752 51484 3758 51536
rect 3142 51456 3148 51468
rect 2884 51428 3148 51456
rect 2409 51391 2467 51397
rect 2409 51357 2421 51391
rect 2455 51357 2467 51391
rect 2409 51351 2467 51357
rect 1688 51292 2268 51320
rect 2424 51320 2452 51351
rect 2774 51348 2780 51400
rect 2832 51388 2838 51400
rect 2884 51397 2912 51428
rect 3142 51416 3148 51428
rect 3200 51416 3206 51468
rect 2869 51391 2927 51397
rect 2869 51388 2881 51391
rect 2832 51360 2881 51388
rect 2832 51348 2838 51360
rect 2869 51357 2881 51360
rect 2915 51357 2927 51391
rect 3050 51388 3056 51400
rect 3011 51360 3056 51388
rect 2869 51351 2927 51357
rect 3050 51348 3056 51360
rect 3108 51348 3114 51400
rect 9858 51388 9864 51400
rect 9819 51360 9864 51388
rect 9858 51348 9864 51360
rect 9916 51348 9922 51400
rect 2958 51320 2964 51332
rect 2424 51292 2964 51320
rect 1688 51264 1716 51292
rect 2958 51280 2964 51292
rect 3016 51280 3022 51332
rect 1394 51212 1400 51264
rect 1452 51252 1458 51264
rect 1489 51255 1547 51261
rect 1489 51252 1501 51255
rect 1452 51224 1501 51252
rect 1452 51212 1458 51224
rect 1489 51221 1501 51224
rect 1535 51221 1547 51255
rect 1489 51215 1547 51221
rect 1670 51212 1676 51264
rect 1728 51212 1734 51264
rect 2222 51252 2228 51264
rect 2183 51224 2228 51252
rect 2222 51212 2228 51224
rect 2280 51212 2286 51264
rect 10042 51252 10048 51264
rect 10003 51224 10048 51252
rect 10042 51212 10048 51224
rect 10100 51212 10106 51264
rect 1104 51162 10856 51184
rect 1104 51110 4213 51162
rect 4265 51110 4277 51162
rect 4329 51110 4341 51162
rect 4393 51110 4405 51162
rect 4457 51110 4469 51162
rect 4521 51110 7477 51162
rect 7529 51110 7541 51162
rect 7593 51110 7605 51162
rect 7657 51110 7669 51162
rect 7721 51110 7733 51162
rect 7785 51110 10856 51162
rect 1104 51088 10856 51110
rect 2222 51008 2228 51060
rect 2280 51048 2286 51060
rect 2869 51051 2927 51057
rect 2280 51020 2325 51048
rect 2280 51008 2286 51020
rect 2869 51017 2881 51051
rect 2915 51048 2927 51051
rect 3234 51048 3240 51060
rect 2915 51020 3240 51048
rect 2915 51017 2927 51020
rect 2869 51011 2927 51017
rect 3234 51008 3240 51020
rect 3292 51008 3298 51060
rect 3694 51048 3700 51060
rect 3436 51020 3700 51048
rect 3050 50980 3056 50992
rect 2608 50952 3056 50980
rect 1673 50915 1731 50921
rect 1673 50881 1685 50915
rect 1719 50881 1731 50915
rect 1673 50875 1731 50881
rect 2133 50915 2191 50921
rect 2133 50881 2145 50915
rect 2179 50912 2191 50915
rect 2222 50912 2228 50924
rect 2179 50884 2228 50912
rect 2179 50881 2191 50884
rect 2133 50875 2191 50881
rect 1688 50844 1716 50875
rect 2222 50872 2228 50884
rect 2280 50872 2286 50924
rect 2317 50915 2375 50921
rect 2317 50881 2329 50915
rect 2363 50912 2375 50915
rect 2498 50912 2504 50924
rect 2363 50884 2504 50912
rect 2363 50881 2375 50884
rect 2317 50875 2375 50881
rect 2498 50872 2504 50884
rect 2556 50872 2562 50924
rect 2608 50844 2636 50952
rect 3050 50940 3056 50952
rect 3108 50940 3114 50992
rect 3436 50980 3464 51020
rect 3694 51008 3700 51020
rect 3752 51008 3758 51060
rect 3160 50952 3464 50980
rect 3513 50983 3571 50989
rect 2774 50912 2780 50924
rect 2735 50884 2780 50912
rect 2774 50872 2780 50884
rect 2832 50872 2838 50924
rect 2961 50915 3019 50921
rect 2961 50881 2973 50915
rect 3007 50912 3019 50915
rect 3160 50912 3188 50952
rect 3513 50949 3525 50983
rect 3559 50980 3571 50983
rect 3559 50952 9904 50980
rect 3559 50949 3571 50952
rect 3513 50943 3571 50949
rect 3421 50915 3479 50921
rect 3421 50912 3433 50915
rect 3007 50884 3188 50912
rect 3252 50884 3433 50912
rect 3007 50881 3019 50884
rect 2961 50875 3019 50881
rect 1688 50816 2636 50844
rect 2792 50844 2820 50872
rect 3050 50844 3056 50856
rect 2792 50816 3056 50844
rect 3050 50804 3056 50816
rect 3108 50804 3114 50856
rect 198 50736 204 50788
rect 256 50776 262 50788
rect 256 50748 1624 50776
rect 256 50736 262 50748
rect 1486 50708 1492 50720
rect 1447 50680 1492 50708
rect 1486 50668 1492 50680
rect 1544 50668 1550 50720
rect 1596 50708 1624 50748
rect 1946 50736 1952 50788
rect 2004 50776 2010 50788
rect 2682 50776 2688 50788
rect 2004 50748 2688 50776
rect 2004 50736 2010 50748
rect 2682 50736 2688 50748
rect 2740 50736 2746 50788
rect 3252 50708 3280 50884
rect 3421 50881 3433 50884
rect 3467 50881 3479 50915
rect 3421 50875 3479 50881
rect 3605 50915 3663 50921
rect 3605 50881 3617 50915
rect 3651 50912 3663 50915
rect 3694 50912 3700 50924
rect 3651 50884 3700 50912
rect 3651 50881 3663 50884
rect 3605 50875 3663 50881
rect 3694 50872 3700 50884
rect 3752 50872 3758 50924
rect 9876 50921 9904 50952
rect 9861 50915 9919 50921
rect 9861 50881 9873 50915
rect 9907 50881 9919 50915
rect 9861 50875 9919 50881
rect 10042 50708 10048 50720
rect 1596 50680 3280 50708
rect 10003 50680 10048 50708
rect 10042 50668 10048 50680
rect 10100 50668 10106 50720
rect 1104 50618 10856 50640
rect 1104 50566 2582 50618
rect 2634 50566 2646 50618
rect 2698 50566 2710 50618
rect 2762 50566 2774 50618
rect 2826 50566 2838 50618
rect 2890 50566 5845 50618
rect 5897 50566 5909 50618
rect 5961 50566 5973 50618
rect 6025 50566 6037 50618
rect 6089 50566 6101 50618
rect 6153 50566 9109 50618
rect 9161 50566 9173 50618
rect 9225 50566 9237 50618
rect 9289 50566 9301 50618
rect 9353 50566 9365 50618
rect 9417 50566 10856 50618
rect 1104 50544 10856 50566
rect 106 50464 112 50516
rect 164 50504 170 50516
rect 1670 50504 1676 50516
rect 164 50476 1676 50504
rect 164 50464 170 50476
rect 1670 50464 1676 50476
rect 1728 50504 1734 50516
rect 3234 50504 3240 50516
rect 1728 50476 3240 50504
rect 1728 50464 1734 50476
rect 3234 50464 3240 50476
rect 3292 50464 3298 50516
rect 3973 50507 4031 50513
rect 3973 50473 3985 50507
rect 4019 50504 4031 50507
rect 4617 50507 4675 50513
rect 4019 50476 4568 50504
rect 4019 50473 4031 50476
rect 3973 50467 4031 50473
rect 1949 50439 2007 50445
rect 1949 50436 1961 50439
rect 1228 50408 1961 50436
rect 1228 50244 1256 50408
rect 1949 50405 1961 50408
rect 1995 50405 2007 50439
rect 1949 50399 2007 50405
rect 2406 50396 2412 50448
rect 2464 50396 2470 50448
rect 4540 50436 4568 50476
rect 4617 50473 4629 50507
rect 4663 50504 4675 50507
rect 9858 50504 9864 50516
rect 4663 50476 9864 50504
rect 4663 50473 4675 50476
rect 4617 50467 4675 50473
rect 9858 50464 9864 50476
rect 9916 50464 9922 50516
rect 10873 50439 10931 50445
rect 4540 50408 9812 50436
rect 1670 50368 1676 50380
rect 1412 50340 1676 50368
rect 1412 50309 1440 50340
rect 1670 50328 1676 50340
rect 1728 50368 1734 50380
rect 2424 50368 2452 50396
rect 1728 50340 2452 50368
rect 2685 50371 2743 50377
rect 1728 50328 1734 50340
rect 2685 50337 2697 50371
rect 2731 50368 2743 50371
rect 3050 50368 3056 50380
rect 2731 50340 3056 50368
rect 2731 50337 2743 50340
rect 2685 50331 2743 50337
rect 3050 50328 3056 50340
rect 3108 50328 3114 50380
rect 1397 50303 1455 50309
rect 1397 50269 1409 50303
rect 1443 50269 1455 50303
rect 1578 50300 1584 50312
rect 1539 50272 1584 50300
rect 1397 50263 1455 50269
rect 1578 50260 1584 50272
rect 1636 50260 1642 50312
rect 1765 50303 1823 50309
rect 1765 50269 1777 50303
rect 1811 50300 1823 50303
rect 1854 50300 1860 50312
rect 1811 50272 1860 50300
rect 1811 50269 1823 50272
rect 1765 50263 1823 50269
rect 1854 50260 1860 50272
rect 1912 50300 1918 50312
rect 2222 50300 2228 50312
rect 1912 50272 2228 50300
rect 1912 50260 1918 50272
rect 2222 50260 2228 50272
rect 2280 50260 2286 50312
rect 2409 50303 2467 50309
rect 2409 50269 2421 50303
rect 2455 50300 2467 50303
rect 2455 50272 3096 50300
rect 2455 50269 2467 50272
rect 2409 50263 2467 50269
rect 3068 50244 3096 50272
rect 3234 50260 3240 50312
rect 3292 50300 3298 50312
rect 3789 50303 3847 50309
rect 3789 50300 3801 50303
rect 3292 50272 3801 50300
rect 3292 50260 3298 50272
rect 3789 50269 3801 50272
rect 3835 50269 3847 50303
rect 3789 50263 3847 50269
rect 3878 50260 3884 50312
rect 3936 50300 3942 50312
rect 3973 50303 4031 50309
rect 3973 50300 3985 50303
rect 3936 50272 3985 50300
rect 3936 50260 3942 50272
rect 3973 50269 3985 50272
rect 4019 50269 4031 50303
rect 3973 50263 4031 50269
rect 4433 50303 4491 50309
rect 4433 50269 4445 50303
rect 4479 50269 4491 50303
rect 4433 50263 4491 50269
rect 4617 50303 4675 50309
rect 4617 50269 4629 50303
rect 4663 50269 4675 50303
rect 4617 50263 4675 50269
rect 1210 50192 1216 50244
rect 1268 50192 1274 50244
rect 1673 50235 1731 50241
rect 1673 50201 1685 50235
rect 1719 50232 1731 50235
rect 2774 50232 2780 50244
rect 1719 50204 2780 50232
rect 1719 50201 1731 50204
rect 1673 50195 1731 50201
rect 2774 50192 2780 50204
rect 2832 50192 2838 50244
rect 3050 50192 3056 50244
rect 3108 50192 3114 50244
rect 3418 50192 3424 50244
rect 3476 50232 3482 50244
rect 4448 50232 4476 50263
rect 3476 50204 4476 50232
rect 3476 50192 3482 50204
rect 937 50167 995 50173
rect 937 50133 949 50167
rect 983 50164 995 50167
rect 1578 50164 1584 50176
rect 983 50136 1584 50164
rect 983 50133 995 50136
rect 937 50127 995 50133
rect 1578 50124 1584 50136
rect 1636 50124 1642 50176
rect 3234 50124 3240 50176
rect 3292 50164 3298 50176
rect 3694 50164 3700 50176
rect 3292 50136 3700 50164
rect 3292 50124 3298 50136
rect 3694 50124 3700 50136
rect 3752 50164 3758 50176
rect 4632 50164 4660 50263
rect 9784 50232 9812 50408
rect 10873 50405 10885 50439
rect 10919 50436 10931 50439
rect 11517 50439 11575 50445
rect 11517 50436 11529 50439
rect 10919 50408 11529 50436
rect 10919 50405 10931 50408
rect 10873 50399 10931 50405
rect 11517 50405 11529 50408
rect 11563 50405 11575 50439
rect 11517 50399 11575 50405
rect 11609 50439 11667 50445
rect 11609 50405 11621 50439
rect 11655 50436 11667 50439
rect 11655 50408 11744 50436
rect 11655 50405 11667 50408
rect 11609 50399 11667 50405
rect 10962 50368 10968 50380
rect 10923 50340 10968 50368
rect 10962 50328 10968 50340
rect 11020 50328 11026 50380
rect 11716 50309 11744 50408
rect 9861 50303 9919 50309
rect 9861 50269 9873 50303
rect 9907 50300 9919 50303
rect 11609 50303 11667 50309
rect 11609 50300 11621 50303
rect 9907 50272 11621 50300
rect 9907 50269 9919 50272
rect 9861 50263 9919 50269
rect 11609 50269 11621 50272
rect 11655 50269 11667 50303
rect 11609 50263 11667 50269
rect 11701 50303 11759 50309
rect 11701 50269 11713 50303
rect 11747 50269 11759 50303
rect 11701 50263 11759 50269
rect 10965 50235 11023 50241
rect 10965 50232 10977 50235
rect 9784 50204 10977 50232
rect 10965 50201 10977 50204
rect 11011 50201 11023 50235
rect 10965 50195 11023 50201
rect 10042 50164 10048 50176
rect 3752 50136 4660 50164
rect 10003 50136 10048 50164
rect 3752 50124 3758 50136
rect 10042 50124 10048 50136
rect 10100 50124 10106 50176
rect 10873 50167 10931 50173
rect 10873 50133 10885 50167
rect 10919 50133 10931 50167
rect 10873 50127 10931 50133
rect 1104 50074 10856 50096
rect 1104 50022 4213 50074
rect 4265 50022 4277 50074
rect 4329 50022 4341 50074
rect 4393 50022 4405 50074
rect 4457 50022 4469 50074
rect 4521 50022 7477 50074
rect 7529 50022 7541 50074
rect 7593 50022 7605 50074
rect 7657 50022 7669 50074
rect 7721 50022 7733 50074
rect 7785 50022 10856 50074
rect 1104 50000 10856 50022
rect 1762 49960 1768 49972
rect 1596 49932 1768 49960
rect 1596 49901 1624 49932
rect 1762 49920 1768 49932
rect 1820 49920 1826 49972
rect 2774 49920 2780 49972
rect 2832 49960 2838 49972
rect 10888 49960 10916 50127
rect 2832 49932 10916 49960
rect 2832 49920 2838 49932
rect 1581 49895 1639 49901
rect 1581 49861 1593 49895
rect 1627 49861 1639 49895
rect 1581 49855 1639 49861
rect 1673 49895 1731 49901
rect 1673 49861 1685 49895
rect 1719 49892 1731 49895
rect 4154 49892 4160 49904
rect 1719 49864 2820 49892
rect 1719 49861 1731 49864
rect 1673 49855 1731 49861
rect 1397 49827 1455 49833
rect 1397 49793 1409 49827
rect 1443 49824 1455 49827
rect 1765 49827 1823 49833
rect 1443 49796 1716 49824
rect 1443 49793 1455 49796
rect 1397 49787 1455 49793
rect 1688 49768 1716 49796
rect 1765 49793 1777 49827
rect 1811 49824 1823 49827
rect 2222 49824 2228 49836
rect 1811 49796 2228 49824
rect 1811 49793 1823 49796
rect 1765 49787 1823 49793
rect 2222 49784 2228 49796
rect 2280 49784 2286 49836
rect 2406 49824 2412 49836
rect 2367 49796 2412 49824
rect 2406 49784 2412 49796
rect 2464 49784 2470 49836
rect 290 49716 296 49768
rect 348 49756 354 49768
rect 348 49728 1624 49756
rect 348 49716 354 49728
rect 1596 49688 1624 49728
rect 1670 49716 1676 49768
rect 1728 49716 1734 49768
rect 1949 49691 2007 49697
rect 1949 49688 1961 49691
rect 1596 49660 1961 49688
rect 1949 49657 1961 49660
rect 1995 49657 2007 49691
rect 1949 49651 2007 49657
rect 2406 49580 2412 49632
rect 2464 49620 2470 49632
rect 2593 49623 2651 49629
rect 2593 49620 2605 49623
rect 2464 49592 2605 49620
rect 2464 49580 2470 49592
rect 2593 49589 2605 49592
rect 2639 49589 2651 49623
rect 2792 49620 2820 49864
rect 3344 49864 4160 49892
rect 3344 49833 3372 49864
rect 4154 49852 4160 49864
rect 4212 49892 4218 49904
rect 4890 49892 4896 49904
rect 4212 49864 4896 49892
rect 4212 49852 4218 49864
rect 4890 49852 4896 49864
rect 4948 49852 4954 49904
rect 3329 49827 3387 49833
rect 3329 49793 3341 49827
rect 3375 49793 3387 49827
rect 3329 49787 3387 49793
rect 3513 49827 3571 49833
rect 3513 49793 3525 49827
rect 3559 49824 3571 49827
rect 3694 49824 3700 49836
rect 3559 49796 3700 49824
rect 3559 49793 3571 49796
rect 3513 49787 3571 49793
rect 3694 49784 3700 49796
rect 3752 49824 3758 49836
rect 3878 49824 3884 49836
rect 3752 49796 3884 49824
rect 3752 49784 3758 49796
rect 3878 49784 3884 49796
rect 3936 49784 3942 49836
rect 6181 49827 6239 49833
rect 6181 49793 6193 49827
rect 6227 49824 6239 49827
rect 10962 49824 10968 49836
rect 6227 49796 10968 49824
rect 6227 49793 6239 49796
rect 6181 49787 6239 49793
rect 10962 49784 10968 49796
rect 11020 49784 11026 49836
rect 3421 49759 3479 49765
rect 3421 49725 3433 49759
rect 3467 49756 3479 49759
rect 9674 49756 9680 49768
rect 3467 49728 4016 49756
rect 3467 49725 3479 49728
rect 3421 49719 3479 49725
rect 3988 49688 4016 49728
rect 9646 49716 9680 49756
rect 9732 49716 9738 49768
rect 9646 49688 9674 49716
rect 3988 49660 9674 49688
rect 6181 49623 6239 49629
rect 6181 49620 6193 49623
rect 2792 49592 6193 49620
rect 2593 49583 2651 49589
rect 6181 49589 6193 49592
rect 6227 49589 6239 49623
rect 6181 49583 6239 49589
rect 11701 49555 11759 49561
rect 11701 49552 11713 49555
rect 1104 49530 10856 49552
rect 1104 49478 2582 49530
rect 2634 49478 2646 49530
rect 2698 49478 2710 49530
rect 2762 49478 2774 49530
rect 2826 49478 2838 49530
rect 2890 49478 5845 49530
rect 5897 49478 5909 49530
rect 5961 49478 5973 49530
rect 6025 49478 6037 49530
rect 6089 49478 6101 49530
rect 6153 49478 9109 49530
rect 9161 49478 9173 49530
rect 9225 49478 9237 49530
rect 9289 49478 9301 49530
rect 9353 49478 9365 49530
rect 9417 49478 10856 49530
rect 1104 49456 10856 49478
rect 10888 49524 11713 49552
rect 658 49376 664 49428
rect 716 49416 722 49428
rect 1578 49416 1584 49428
rect 716 49388 1584 49416
rect 716 49376 722 49388
rect 1578 49376 1584 49388
rect 1636 49376 1642 49428
rect 1762 49376 1768 49428
rect 1820 49416 1826 49428
rect 1946 49416 1952 49428
rect 1820 49388 1952 49416
rect 1820 49376 1826 49388
rect 1946 49376 1952 49388
rect 2004 49376 2010 49428
rect 4798 49376 4804 49428
rect 4856 49416 4862 49428
rect 5166 49416 5172 49428
rect 4856 49388 5172 49416
rect 4856 49376 4862 49388
rect 5166 49376 5172 49388
rect 5224 49376 5230 49428
rect 2222 49348 2228 49360
rect 1596 49320 2228 49348
rect 1394 49172 1400 49224
rect 1452 49172 1458 49224
rect 1596 49221 1624 49320
rect 2222 49308 2228 49320
rect 2280 49308 2286 49360
rect 10888 49348 10916 49524
rect 11701 49521 11713 49524
rect 11747 49521 11759 49555
rect 11701 49515 11759 49521
rect 11149 49419 11207 49425
rect 11149 49385 11161 49419
rect 11195 49416 11207 49419
rect 11701 49419 11759 49425
rect 11701 49416 11713 49419
rect 11195 49388 11713 49416
rect 11195 49385 11207 49388
rect 11149 49379 11207 49385
rect 11701 49385 11713 49388
rect 11747 49385 11759 49419
rect 11701 49379 11759 49385
rect 2746 49320 10916 49348
rect 2746 49280 2774 49320
rect 3878 49280 3884 49292
rect 1688 49252 2774 49280
rect 3791 49252 3884 49280
rect 1688 49221 1716 49252
rect 1581 49215 1639 49221
rect 1581 49181 1593 49215
rect 1627 49181 1639 49215
rect 1581 49175 1639 49181
rect 1673 49215 1731 49221
rect 1673 49181 1685 49215
rect 1719 49181 1731 49215
rect 1946 49212 1952 49224
rect 1907 49184 1952 49212
rect 1673 49175 1731 49181
rect 1946 49172 1952 49184
rect 2004 49172 2010 49224
rect 2682 49212 2688 49224
rect 2643 49184 2688 49212
rect 2682 49172 2688 49184
rect 2740 49172 2746 49224
rect 3804 49221 3832 49252
rect 3878 49240 3884 49252
rect 3936 49280 3942 49292
rect 5166 49280 5172 49292
rect 3936 49252 5172 49280
rect 3936 49240 3942 49252
rect 5166 49240 5172 49252
rect 5224 49240 5230 49292
rect 3789 49215 3847 49221
rect 3789 49181 3801 49215
rect 3835 49181 3847 49215
rect 3789 49175 3847 49181
rect 3973 49215 4031 49221
rect 3973 49181 3985 49215
rect 4019 49181 4031 49215
rect 3973 49175 4031 49181
rect 1412 49144 1440 49172
rect 1765 49147 1823 49153
rect 1765 49144 1777 49147
rect 1412 49116 1777 49144
rect 1765 49113 1777 49116
rect 1811 49113 1823 49147
rect 1765 49107 1823 49113
rect 3694 49104 3700 49156
rect 3752 49144 3758 49156
rect 3988 49144 4016 49175
rect 9582 49172 9588 49224
rect 9640 49212 9646 49224
rect 9861 49215 9919 49221
rect 9861 49212 9873 49215
rect 9640 49184 9873 49212
rect 9640 49172 9646 49184
rect 9861 49181 9873 49184
rect 9907 49181 9919 49215
rect 9861 49175 9919 49181
rect 3752 49116 4016 49144
rect 3752 49104 3758 49116
rect 1394 49076 1400 49088
rect 1355 49048 1400 49076
rect 1394 49036 1400 49048
rect 1452 49036 1458 49088
rect 2501 49079 2559 49085
rect 2501 49045 2513 49079
rect 2547 49076 2559 49079
rect 2774 49076 2780 49088
rect 2547 49048 2780 49076
rect 2547 49045 2559 49048
rect 2501 49039 2559 49045
rect 2774 49036 2780 49048
rect 2832 49036 2838 49088
rect 3881 49079 3939 49085
rect 3881 49045 3893 49079
rect 3927 49076 3939 49079
rect 9858 49076 9864 49088
rect 3927 49048 9864 49076
rect 3927 49045 3939 49048
rect 3881 49039 3939 49045
rect 9858 49036 9864 49048
rect 9916 49036 9922 49088
rect 10042 49076 10048 49088
rect 10003 49048 10048 49076
rect 10042 49036 10048 49048
rect 10100 49036 10106 49088
rect 1104 48986 10856 49008
rect 1104 48934 4213 48986
rect 4265 48934 4277 48986
rect 4329 48934 4341 48986
rect 4393 48934 4405 48986
rect 4457 48934 4469 48986
rect 4521 48934 7477 48986
rect 7529 48934 7541 48986
rect 7593 48934 7605 48986
rect 7657 48934 7669 48986
rect 7721 48934 7733 48986
rect 7785 48934 10856 48986
rect 1104 48912 10856 48934
rect 2222 48872 2228 48884
rect 2183 48844 2228 48872
rect 2222 48832 2228 48844
rect 2280 48832 2286 48884
rect 2682 48832 2688 48884
rect 2740 48872 2746 48884
rect 6454 48872 6460 48884
rect 2740 48844 6460 48872
rect 2740 48832 2746 48844
rect 6454 48832 6460 48844
rect 6512 48832 6518 48884
rect 658 48764 664 48816
rect 716 48804 722 48816
rect 1946 48804 1952 48816
rect 716 48776 1952 48804
rect 716 48764 722 48776
rect 1946 48764 1952 48776
rect 2004 48804 2010 48816
rect 2004 48776 3280 48804
rect 2004 48764 2010 48776
rect 1673 48739 1731 48745
rect 1673 48705 1685 48739
rect 1719 48736 1731 48739
rect 2222 48736 2228 48748
rect 1719 48708 2228 48736
rect 1719 48705 1731 48708
rect 1673 48699 1731 48705
rect 2222 48696 2228 48708
rect 2280 48696 2286 48748
rect 3252 48745 3280 48776
rect 2409 48739 2467 48745
rect 2409 48705 2421 48739
rect 2455 48705 2467 48739
rect 2409 48699 2467 48705
rect 3237 48739 3295 48745
rect 3237 48705 3249 48739
rect 3283 48705 3295 48739
rect 3237 48699 3295 48705
rect 3421 48739 3479 48745
rect 3421 48705 3433 48739
rect 3467 48736 3479 48739
rect 3694 48736 3700 48748
rect 3467 48708 3700 48736
rect 3467 48705 3479 48708
rect 3421 48699 3479 48705
rect 1486 48532 1492 48544
rect 1447 48504 1492 48532
rect 1486 48492 1492 48504
rect 1544 48492 1550 48544
rect 2424 48532 2452 48699
rect 3694 48696 3700 48708
rect 3752 48696 3758 48748
rect 9766 48696 9772 48748
rect 9824 48736 9830 48748
rect 9861 48739 9919 48745
rect 9861 48736 9873 48739
rect 9824 48708 9873 48736
rect 9824 48696 9830 48708
rect 9861 48705 9873 48708
rect 9907 48705 9919 48739
rect 9861 48699 9919 48705
rect 3329 48671 3387 48677
rect 3329 48637 3341 48671
rect 3375 48668 3387 48671
rect 3375 48640 6224 48668
rect 3375 48637 3387 48640
rect 3329 48631 3387 48637
rect 6086 48560 6092 48612
rect 6144 48560 6150 48612
rect 6196 48600 6224 48640
rect 10965 48603 11023 48609
rect 10965 48600 10977 48603
rect 6196 48572 6316 48600
rect 5718 48532 5724 48544
rect 2424 48504 5724 48532
rect 5718 48492 5724 48504
rect 5776 48492 5782 48544
rect 6104 48532 6132 48560
rect 6178 48532 6184 48544
rect 6104 48504 6184 48532
rect 6178 48492 6184 48504
rect 6236 48492 6242 48544
rect 6288 48532 6316 48572
rect 9646 48572 10977 48600
rect 9646 48532 9674 48572
rect 10965 48569 10977 48572
rect 11011 48569 11023 48603
rect 10965 48563 11023 48569
rect 10042 48532 10048 48544
rect 6288 48504 9674 48532
rect 10003 48504 10048 48532
rect 10042 48492 10048 48504
rect 10100 48492 10106 48544
rect 1104 48442 10856 48464
rect 1104 48390 2582 48442
rect 2634 48390 2646 48442
rect 2698 48390 2710 48442
rect 2762 48390 2774 48442
rect 2826 48390 2838 48442
rect 2890 48390 5845 48442
rect 5897 48390 5909 48442
rect 5961 48390 5973 48442
rect 6025 48390 6037 48442
rect 6089 48390 6101 48442
rect 6153 48390 9109 48442
rect 9161 48390 9173 48442
rect 9225 48390 9237 48442
rect 9289 48390 9301 48442
rect 9353 48390 9365 48442
rect 9417 48390 10856 48442
rect 1104 48368 10856 48390
rect 382 48288 388 48340
rect 440 48328 446 48340
rect 2406 48328 2412 48340
rect 440 48300 2412 48328
rect 440 48288 446 48300
rect 2406 48288 2412 48300
rect 2464 48288 2470 48340
rect 4614 48328 4620 48340
rect 2700 48300 4620 48328
rect 2700 48272 2728 48300
rect 4614 48288 4620 48300
rect 4672 48288 4678 48340
rect 2682 48220 2688 48272
rect 2740 48220 2746 48272
rect 2961 48263 3019 48269
rect 2961 48229 2973 48263
rect 3007 48260 3019 48263
rect 9766 48260 9772 48272
rect 3007 48232 5580 48260
rect 3007 48229 3019 48232
rect 2961 48223 3019 48229
rect 198 48152 204 48204
rect 256 48192 262 48204
rect 2225 48195 2283 48201
rect 256 48164 2176 48192
rect 256 48152 262 48164
rect 1673 48127 1731 48133
rect 1673 48093 1685 48127
rect 1719 48124 1731 48127
rect 2038 48124 2044 48136
rect 1719 48096 2044 48124
rect 1719 48093 1731 48096
rect 1673 48087 1731 48093
rect 2038 48084 2044 48096
rect 2096 48084 2102 48136
rect 2148 48133 2176 48164
rect 2225 48161 2237 48195
rect 2271 48192 2283 48195
rect 5074 48192 5080 48204
rect 2271 48164 5080 48192
rect 2271 48161 2283 48164
rect 2225 48155 2283 48161
rect 5074 48152 5080 48164
rect 5132 48152 5138 48204
rect 5552 48192 5580 48232
rect 8266 48232 9772 48260
rect 8266 48192 8294 48232
rect 9766 48220 9772 48232
rect 9824 48220 9830 48272
rect 5552 48164 8294 48192
rect 2133 48127 2191 48133
rect 2133 48093 2145 48127
rect 2179 48093 2191 48127
rect 2133 48087 2191 48093
rect 2317 48127 2375 48133
rect 2317 48093 2329 48127
rect 2363 48093 2375 48127
rect 2317 48087 2375 48093
rect 2777 48127 2835 48133
rect 2777 48093 2789 48127
rect 2823 48093 2835 48127
rect 2777 48087 2835 48093
rect 2961 48127 3019 48133
rect 2961 48093 2973 48127
rect 3007 48124 3019 48127
rect 3234 48124 3240 48136
rect 3007 48096 3240 48124
rect 3007 48093 3019 48096
rect 2961 48087 3019 48093
rect 382 48016 388 48068
rect 440 48056 446 48068
rect 440 48028 1624 48056
rect 440 48016 446 48028
rect 1486 47988 1492 48000
rect 1447 47960 1492 47988
rect 1486 47948 1492 47960
rect 1544 47948 1550 48000
rect 1596 47988 1624 48028
rect 1762 48016 1768 48068
rect 1820 48056 1826 48068
rect 2332 48056 2360 48087
rect 1820 48028 2360 48056
rect 1820 48016 1826 48028
rect 2792 47988 2820 48087
rect 3234 48084 3240 48096
rect 3292 48084 3298 48136
rect 3142 47988 3148 48000
rect 1596 47960 3148 47988
rect 3142 47948 3148 47960
rect 3200 47948 3206 48000
rect 1104 47898 10856 47920
rect 1104 47846 4213 47898
rect 4265 47846 4277 47898
rect 4329 47846 4341 47898
rect 4393 47846 4405 47898
rect 4457 47846 4469 47898
rect 4521 47846 7477 47898
rect 7529 47846 7541 47898
rect 7593 47846 7605 47898
rect 7657 47846 7669 47898
rect 7721 47846 7733 47898
rect 7785 47846 10856 47898
rect 1104 47824 10856 47846
rect 2869 47787 2927 47793
rect 2869 47753 2881 47787
rect 2915 47784 2927 47787
rect 2958 47784 2964 47796
rect 2915 47756 2964 47784
rect 2915 47753 2927 47756
rect 2869 47747 2927 47753
rect 2958 47744 2964 47756
rect 3016 47744 3022 47796
rect 2038 47676 2044 47728
rect 2096 47716 2102 47728
rect 6178 47716 6184 47728
rect 2096 47688 6184 47716
rect 2096 47676 2102 47688
rect 6178 47676 6184 47688
rect 6236 47676 6242 47728
rect 1673 47651 1731 47657
rect 1673 47617 1685 47651
rect 1719 47617 1731 47651
rect 1673 47611 1731 47617
rect 2409 47651 2467 47657
rect 2409 47617 2421 47651
rect 2455 47648 2467 47651
rect 3053 47651 3111 47657
rect 2455 47620 2774 47648
rect 2455 47617 2467 47620
rect 2409 47611 2467 47617
rect 1688 47512 1716 47611
rect 2746 47580 2774 47620
rect 3053 47617 3065 47651
rect 3099 47648 3111 47651
rect 3142 47648 3148 47660
rect 3099 47620 3148 47648
rect 3099 47617 3111 47620
rect 3053 47611 3111 47617
rect 3142 47608 3148 47620
rect 3200 47608 3206 47660
rect 9674 47608 9680 47660
rect 9732 47648 9738 47660
rect 9861 47651 9919 47657
rect 9861 47648 9873 47651
rect 9732 47620 9873 47648
rect 9732 47608 9738 47620
rect 9861 47617 9873 47620
rect 9907 47617 9919 47651
rect 9861 47611 9919 47617
rect 7926 47580 7932 47592
rect 2746 47552 7932 47580
rect 7926 47540 7932 47552
rect 7984 47540 7990 47592
rect 9030 47512 9036 47524
rect 1688 47484 9036 47512
rect 9030 47472 9036 47484
rect 9088 47472 9094 47524
rect 10042 47512 10048 47524
rect 10003 47484 10048 47512
rect 10042 47472 10048 47484
rect 10100 47472 10106 47524
rect 1486 47444 1492 47456
rect 1447 47416 1492 47444
rect 1486 47404 1492 47416
rect 1544 47404 1550 47456
rect 2222 47444 2228 47456
rect 2183 47416 2228 47444
rect 2222 47404 2228 47416
rect 2280 47404 2286 47456
rect 1104 47354 10856 47376
rect 1104 47302 2582 47354
rect 2634 47302 2646 47354
rect 2698 47302 2710 47354
rect 2762 47302 2774 47354
rect 2826 47302 2838 47354
rect 2890 47302 5845 47354
rect 5897 47302 5909 47354
rect 5961 47302 5973 47354
rect 6025 47302 6037 47354
rect 6089 47302 6101 47354
rect 6153 47302 9109 47354
rect 9161 47302 9173 47354
rect 9225 47302 9237 47354
rect 9289 47302 9301 47354
rect 9353 47302 9365 47354
rect 9417 47302 10856 47354
rect 1104 47280 10856 47302
rect 2133 47243 2191 47249
rect 2133 47209 2145 47243
rect 2179 47240 2191 47243
rect 2314 47240 2320 47252
rect 2179 47212 2320 47240
rect 2179 47209 2191 47212
rect 2133 47203 2191 47209
rect 2314 47200 2320 47212
rect 2372 47200 2378 47252
rect 2961 47243 3019 47249
rect 2961 47209 2973 47243
rect 3007 47240 3019 47243
rect 3786 47240 3792 47252
rect 3007 47212 3792 47240
rect 3007 47209 3019 47212
rect 2961 47203 3019 47209
rect 3786 47200 3792 47212
rect 3844 47200 3850 47252
rect 4614 47132 4620 47184
rect 4672 47172 4678 47184
rect 4798 47172 4804 47184
rect 4672 47144 4804 47172
rect 4672 47132 4678 47144
rect 4798 47132 4804 47144
rect 4856 47132 4862 47184
rect 8938 47104 8944 47116
rect 1688 47076 8944 47104
rect 1688 47045 1716 47076
rect 8938 47064 8944 47076
rect 8996 47064 9002 47116
rect 1673 47039 1731 47045
rect 1673 47005 1685 47039
rect 1719 47005 1731 47039
rect 1673 46999 1731 47005
rect 2133 47039 2191 47045
rect 2133 47005 2145 47039
rect 2179 47005 2191 47039
rect 2314 47036 2320 47048
rect 2275 47008 2320 47036
rect 2133 46999 2191 47005
rect 2148 46968 2176 46999
rect 2314 46996 2320 47008
rect 2372 46996 2378 47048
rect 2961 47039 3019 47045
rect 2961 47005 2973 47039
rect 3007 47036 3019 47039
rect 4798 47036 4804 47048
rect 3007 47008 4804 47036
rect 3007 47005 3019 47008
rect 2961 46999 3019 47005
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 9861 47039 9919 47045
rect 9861 47005 9873 47039
rect 9907 47036 9919 47039
rect 11057 47039 11115 47045
rect 11057 47036 11069 47039
rect 9907 47008 11069 47036
rect 9907 47005 9919 47008
rect 9861 46999 9919 47005
rect 11057 47005 11069 47008
rect 11103 47005 11115 47039
rect 11057 46999 11115 47005
rect 2148 46940 2452 46968
rect 1486 46900 1492 46912
rect 1447 46872 1492 46900
rect 1486 46860 1492 46872
rect 1544 46860 1550 46912
rect 2424 46900 2452 46940
rect 2958 46900 2964 46912
rect 2424 46872 2964 46900
rect 2958 46860 2964 46872
rect 3016 46860 3022 46912
rect 10042 46900 10048 46912
rect 10003 46872 10048 46900
rect 10042 46860 10048 46872
rect 10100 46860 10106 46912
rect 1104 46810 10856 46832
rect 1104 46758 4213 46810
rect 4265 46758 4277 46810
rect 4329 46758 4341 46810
rect 4393 46758 4405 46810
rect 4457 46758 4469 46810
rect 4521 46758 7477 46810
rect 7529 46758 7541 46810
rect 7593 46758 7605 46810
rect 7657 46758 7669 46810
rect 7721 46758 7733 46810
rect 7785 46758 10856 46810
rect 1104 46736 10856 46758
rect 1946 46656 1952 46708
rect 2004 46696 2010 46708
rect 2317 46699 2375 46705
rect 2317 46696 2329 46699
rect 2004 46668 2329 46696
rect 2004 46656 2010 46668
rect 2317 46665 2329 46668
rect 2363 46665 2375 46699
rect 2317 46659 2375 46665
rect 2406 46656 2412 46708
rect 2464 46696 2470 46708
rect 2590 46696 2596 46708
rect 2464 46668 2596 46696
rect 2464 46656 2470 46668
rect 2590 46656 2596 46668
rect 2648 46656 2654 46708
rect 2961 46699 3019 46705
rect 2961 46665 2973 46699
rect 3007 46696 3019 46699
rect 9582 46696 9588 46708
rect 3007 46668 9588 46696
rect 3007 46665 3019 46668
rect 2961 46659 3019 46665
rect 9582 46656 9588 46668
rect 9640 46656 9646 46708
rect 1673 46563 1731 46569
rect 1673 46529 1685 46563
rect 1719 46529 1731 46563
rect 1673 46523 1731 46529
rect 2225 46563 2283 46569
rect 2225 46529 2237 46563
rect 2271 46529 2283 46563
rect 2225 46523 2283 46529
rect 2409 46563 2467 46569
rect 2409 46529 2421 46563
rect 2455 46529 2467 46563
rect 2409 46523 2467 46529
rect 1486 46356 1492 46368
rect 1447 46328 1492 46356
rect 1486 46316 1492 46328
rect 1544 46316 1550 46368
rect 1688 46356 1716 46523
rect 2240 46424 2268 46523
rect 2424 46492 2452 46523
rect 2590 46520 2596 46572
rect 2648 46560 2654 46572
rect 2869 46563 2927 46569
rect 2869 46560 2881 46563
rect 2648 46532 2881 46560
rect 2648 46520 2654 46532
rect 2869 46529 2881 46532
rect 2915 46529 2927 46563
rect 2869 46523 2927 46529
rect 2958 46520 2964 46572
rect 3016 46520 3022 46572
rect 3053 46563 3111 46569
rect 3053 46529 3065 46563
rect 3099 46560 3111 46563
rect 3234 46560 3240 46572
rect 3099 46532 3240 46560
rect 3099 46529 3111 46532
rect 3053 46523 3111 46529
rect 3234 46520 3240 46532
rect 3292 46560 3298 46572
rect 3878 46560 3884 46572
rect 3292 46532 3884 46560
rect 3292 46520 3298 46532
rect 3878 46520 3884 46532
rect 3936 46520 3942 46572
rect 9858 46560 9864 46572
rect 9819 46532 9864 46560
rect 9858 46520 9864 46532
rect 9916 46520 9922 46572
rect 2976 46492 3004 46520
rect 2424 46464 3004 46492
rect 3234 46424 3240 46436
rect 2240 46396 3240 46424
rect 3234 46384 3240 46396
rect 3292 46384 3298 46436
rect 4706 46384 4712 46436
rect 4764 46424 4770 46436
rect 5166 46424 5172 46436
rect 4764 46396 5172 46424
rect 4764 46384 4770 46396
rect 5166 46384 5172 46396
rect 5224 46384 5230 46436
rect 4614 46356 4620 46368
rect 1688 46328 4620 46356
rect 4614 46316 4620 46328
rect 4672 46316 4678 46368
rect 10042 46356 10048 46368
rect 10003 46328 10048 46356
rect 10042 46316 10048 46328
rect 10100 46316 10106 46368
rect 11057 46359 11115 46365
rect 11057 46325 11069 46359
rect 11103 46356 11115 46359
rect 11517 46359 11575 46365
rect 11517 46356 11529 46359
rect 11103 46328 11529 46356
rect 11103 46325 11115 46328
rect 11057 46319 11115 46325
rect 11517 46325 11529 46328
rect 11563 46325 11575 46359
rect 11517 46319 11575 46325
rect 1104 46266 10856 46288
rect 1104 46214 2582 46266
rect 2634 46214 2646 46266
rect 2698 46214 2710 46266
rect 2762 46214 2774 46266
rect 2826 46214 2838 46266
rect 2890 46214 5845 46266
rect 5897 46214 5909 46266
rect 5961 46214 5973 46266
rect 6025 46214 6037 46266
rect 6089 46214 6101 46266
rect 6153 46214 9109 46266
rect 9161 46214 9173 46266
rect 9225 46214 9237 46266
rect 9289 46214 9301 46266
rect 9353 46214 9365 46266
rect 9417 46214 10856 46266
rect 1104 46192 10856 46214
rect 11517 46223 11575 46229
rect 11517 46189 11529 46223
rect 11563 46220 11575 46223
rect 11885 46223 11943 46229
rect 11885 46220 11897 46223
rect 11563 46192 11897 46220
rect 11563 46189 11575 46192
rect 11517 46183 11575 46189
rect 11885 46189 11897 46192
rect 11931 46189 11943 46223
rect 11885 46183 11943 46189
rect 1854 46112 1860 46164
rect 1912 46152 1918 46164
rect 2130 46152 2136 46164
rect 1912 46124 2136 46152
rect 1912 46112 1918 46124
rect 2130 46112 2136 46124
rect 2188 46112 2194 46164
rect 7834 46152 7840 46164
rect 7116 46124 7840 46152
rect 4706 46044 4712 46096
rect 4764 46084 4770 46096
rect 5258 46084 5264 46096
rect 4764 46056 5264 46084
rect 4764 46044 4770 46056
rect 5258 46044 5264 46056
rect 5316 46044 5322 46096
rect 5718 46044 5724 46096
rect 5776 46084 5782 46096
rect 6638 46084 6644 46096
rect 5776 46056 6644 46084
rect 5776 46044 5782 46056
rect 6638 46044 6644 46056
rect 6696 46044 6702 46096
rect 474 45976 480 46028
rect 532 46016 538 46028
rect 1673 46019 1731 46025
rect 1673 46016 1685 46019
rect 532 45988 1685 46016
rect 532 45976 538 45988
rect 1673 45985 1685 45988
rect 1719 45985 1731 46019
rect 1673 45979 1731 45985
rect 4890 45976 4896 46028
rect 4948 46016 4954 46028
rect 5442 46016 5448 46028
rect 4948 45988 5448 46016
rect 4948 45976 4954 45988
rect 5442 45976 5448 45988
rect 5500 45976 5506 46028
rect 1762 45948 1768 45960
rect 1723 45920 1768 45948
rect 1762 45908 1768 45920
rect 1820 45908 1826 45960
rect 2041 45951 2099 45957
rect 2041 45917 2053 45951
rect 2087 45948 2099 45951
rect 2130 45948 2136 45960
rect 2087 45920 2136 45948
rect 2087 45917 2099 45920
rect 2041 45911 2099 45917
rect 2130 45908 2136 45920
rect 2188 45908 2194 45960
rect 2314 45908 2320 45960
rect 2372 45948 2378 45960
rect 2501 45951 2559 45957
rect 2501 45948 2513 45951
rect 2372 45920 2513 45948
rect 2372 45908 2378 45920
rect 2501 45917 2513 45920
rect 2547 45917 2559 45951
rect 2501 45911 2559 45917
rect 4522 45840 4528 45892
rect 4580 45880 4586 45892
rect 5442 45880 5448 45892
rect 4580 45852 5448 45880
rect 4580 45840 4586 45852
rect 5442 45840 5448 45852
rect 5500 45840 5506 45892
rect 7116 45824 7144 46124
rect 7834 46112 7840 46124
rect 7892 46112 7898 46164
rect 7282 46084 7288 46096
rect 7208 46056 7288 46084
rect 7208 45824 7236 46056
rect 7282 46044 7288 46056
rect 7340 46044 7346 46096
rect 7374 46044 7380 46096
rect 7432 46084 7438 46096
rect 7926 46084 7932 46096
rect 7432 46056 7932 46084
rect 7432 46044 7438 46056
rect 7926 46044 7932 46056
rect 7984 46044 7990 46096
rect 1946 45772 1952 45824
rect 2004 45812 2010 45824
rect 2406 45812 2412 45824
rect 2004 45784 2412 45812
rect 2004 45772 2010 45784
rect 2406 45772 2412 45784
rect 2464 45772 2470 45824
rect 2685 45815 2743 45821
rect 2685 45781 2697 45815
rect 2731 45812 2743 45815
rect 2958 45812 2964 45824
rect 2731 45784 2964 45812
rect 2731 45781 2743 45784
rect 2685 45775 2743 45781
rect 2958 45772 2964 45784
rect 3016 45772 3022 45824
rect 7098 45772 7104 45824
rect 7156 45772 7162 45824
rect 7190 45772 7196 45824
rect 7248 45772 7254 45824
rect 1104 45722 10856 45744
rect 1104 45670 4213 45722
rect 4265 45670 4277 45722
rect 4329 45670 4341 45722
rect 4393 45670 4405 45722
rect 4457 45670 4469 45722
rect 4521 45670 7477 45722
rect 7529 45670 7541 45722
rect 7593 45670 7605 45722
rect 7657 45670 7669 45722
rect 7721 45670 7733 45722
rect 7785 45670 10856 45722
rect 1104 45648 10856 45670
rect 1673 45475 1731 45481
rect 1673 45441 1685 45475
rect 1719 45472 1731 45475
rect 7926 45472 7932 45484
rect 1719 45444 7932 45472
rect 1719 45441 1731 45444
rect 1673 45435 1731 45441
rect 7926 45432 7932 45444
rect 7984 45432 7990 45484
rect 9861 45475 9919 45481
rect 9861 45441 9873 45475
rect 9907 45472 9919 45475
rect 10965 45475 11023 45481
rect 10965 45472 10977 45475
rect 9907 45444 10977 45472
rect 9907 45441 9919 45444
rect 9861 45435 9919 45441
rect 10965 45441 10977 45444
rect 11011 45441 11023 45475
rect 10965 45435 11023 45441
rect 3418 45404 3424 45416
rect 3379 45376 3424 45404
rect 3418 45364 3424 45376
rect 3476 45364 3482 45416
rect 3694 45404 3700 45416
rect 3655 45376 3700 45404
rect 3694 45364 3700 45376
rect 3752 45364 3758 45416
rect 1486 45268 1492 45280
rect 1447 45240 1492 45268
rect 1486 45228 1492 45240
rect 1544 45228 1550 45280
rect 10042 45268 10048 45280
rect 10003 45240 10048 45268
rect 10042 45228 10048 45240
rect 10100 45228 10106 45280
rect 1104 45178 10856 45200
rect 1104 45126 2582 45178
rect 2634 45126 2646 45178
rect 2698 45126 2710 45178
rect 2762 45126 2774 45178
rect 2826 45126 2838 45178
rect 2890 45126 5845 45178
rect 5897 45126 5909 45178
rect 5961 45126 5973 45178
rect 6025 45126 6037 45178
rect 6089 45126 6101 45178
rect 6153 45126 9109 45178
rect 9161 45126 9173 45178
rect 9225 45126 9237 45178
rect 9289 45126 9301 45178
rect 9353 45126 9365 45178
rect 9417 45126 10856 45178
rect 1104 45104 10856 45126
rect 1026 44888 1032 44940
rect 1084 44928 1090 44940
rect 1489 44931 1547 44937
rect 1489 44928 1501 44931
rect 1084 44900 1501 44928
rect 1084 44888 1090 44900
rect 1489 44897 1501 44900
rect 1535 44897 1547 44931
rect 2038 44928 2044 44940
rect 1489 44891 1547 44897
rect 1872 44900 2044 44928
rect 1673 44863 1731 44869
rect 1673 44829 1685 44863
rect 1719 44860 1731 44863
rect 1762 44860 1768 44872
rect 1719 44832 1768 44860
rect 1719 44829 1731 44832
rect 1673 44823 1731 44829
rect 1762 44820 1768 44832
rect 1820 44820 1826 44872
rect 1872 44869 1900 44900
rect 2038 44888 2044 44900
rect 2096 44928 2102 44940
rect 2406 44928 2412 44940
rect 2096 44900 2412 44928
rect 2096 44888 2102 44900
rect 2406 44888 2412 44900
rect 2464 44888 2470 44940
rect 1857 44863 1915 44869
rect 1857 44829 1869 44863
rect 1903 44829 1915 44863
rect 1857 44823 1915 44829
rect 2593 44863 2651 44869
rect 2593 44829 2605 44863
rect 2639 44860 2651 44863
rect 2958 44860 2964 44872
rect 2639 44832 2964 44860
rect 2639 44829 2651 44832
rect 2593 44823 2651 44829
rect 2958 44820 2964 44832
rect 3016 44820 3022 44872
rect 3053 44863 3111 44869
rect 3053 44829 3065 44863
rect 3099 44829 3111 44863
rect 3053 44823 3111 44829
rect 3237 44863 3295 44869
rect 3237 44829 3249 44863
rect 3283 44860 3295 44863
rect 3694 44860 3700 44872
rect 3283 44832 3700 44860
rect 3283 44829 3295 44832
rect 3237 44823 3295 44829
rect 2406 44724 2412 44736
rect 2367 44696 2412 44724
rect 2406 44684 2412 44696
rect 2464 44684 2470 44736
rect 3068 44724 3096 44823
rect 3694 44820 3700 44832
rect 3752 44820 3758 44872
rect 3786 44820 3792 44872
rect 3844 44860 3850 44872
rect 3973 44863 4031 44869
rect 3844 44832 3889 44860
rect 3844 44820 3850 44832
rect 3973 44829 3985 44863
rect 4019 44860 4031 44863
rect 5074 44860 5080 44872
rect 4019 44832 5080 44860
rect 4019 44829 4031 44832
rect 3973 44823 4031 44829
rect 5074 44820 5080 44832
rect 5132 44820 5138 44872
rect 9861 44863 9919 44869
rect 9861 44829 9873 44863
rect 9907 44829 9919 44863
rect 9861 44823 9919 44829
rect 3145 44795 3203 44801
rect 3145 44761 3157 44795
rect 3191 44792 3203 44795
rect 9876 44792 9904 44823
rect 3191 44764 9904 44792
rect 3191 44761 3203 44764
rect 3145 44755 3203 44761
rect 3234 44724 3240 44736
rect 3068 44696 3240 44724
rect 3234 44684 3240 44696
rect 3292 44724 3298 44736
rect 3694 44724 3700 44736
rect 3292 44696 3700 44724
rect 3292 44684 3298 44696
rect 3694 44684 3700 44696
rect 3752 44684 3758 44736
rect 3881 44727 3939 44733
rect 3881 44693 3893 44727
rect 3927 44724 3939 44727
rect 9858 44724 9864 44736
rect 3927 44696 9864 44724
rect 3927 44693 3939 44696
rect 3881 44687 3939 44693
rect 9858 44684 9864 44696
rect 9916 44684 9922 44736
rect 10042 44724 10048 44736
rect 10003 44696 10048 44724
rect 10042 44684 10048 44696
rect 10100 44684 10106 44736
rect 1104 44634 10856 44656
rect 1104 44582 4213 44634
rect 4265 44582 4277 44634
rect 4329 44582 4341 44634
rect 4393 44582 4405 44634
rect 4457 44582 4469 44634
rect 4521 44582 7477 44634
rect 7529 44582 7541 44634
rect 7593 44582 7605 44634
rect 7657 44582 7669 44634
rect 7721 44582 7733 44634
rect 7785 44582 10856 44634
rect 1104 44560 10856 44582
rect 1118 44480 1124 44532
rect 1176 44520 1182 44532
rect 3145 44523 3203 44529
rect 1176 44492 2360 44520
rect 1176 44480 1182 44492
rect 1504 44424 2268 44452
rect 1504 44393 1532 44424
rect 845 44387 903 44393
rect 845 44353 857 44387
rect 891 44384 903 44387
rect 1489 44387 1547 44393
rect 1489 44384 1501 44387
rect 891 44356 1501 44384
rect 891 44353 903 44356
rect 845 44347 903 44353
rect 1489 44353 1501 44356
rect 1535 44353 1547 44387
rect 1489 44347 1547 44353
rect 1673 44387 1731 44393
rect 1673 44353 1685 44387
rect 1719 44384 1731 44387
rect 1762 44384 1768 44396
rect 1719 44356 1768 44384
rect 1719 44353 1731 44356
rect 1673 44347 1731 44353
rect 937 44251 995 44257
rect 937 44217 949 44251
rect 983 44248 995 44251
rect 1688 44248 1716 44347
rect 1762 44344 1768 44356
rect 1820 44344 1826 44396
rect 2240 44316 2268 44424
rect 2332 44393 2360 44492
rect 3145 44489 3157 44523
rect 3191 44520 3203 44523
rect 3326 44520 3332 44532
rect 3191 44492 3332 44520
rect 3191 44489 3203 44492
rect 3145 44483 3203 44489
rect 3326 44480 3332 44492
rect 3384 44480 3390 44532
rect 3602 44480 3608 44532
rect 3660 44520 3666 44532
rect 3789 44523 3847 44529
rect 3789 44520 3801 44523
rect 3660 44492 3801 44520
rect 3660 44480 3666 44492
rect 3789 44489 3801 44492
rect 3835 44489 3847 44523
rect 3789 44483 3847 44489
rect 4433 44523 4491 44529
rect 4433 44489 4445 44523
rect 4479 44520 4491 44523
rect 11609 44523 11667 44529
rect 11609 44520 11621 44523
rect 4479 44492 11621 44520
rect 4479 44489 4491 44492
rect 4433 44483 4491 44489
rect 11609 44489 11621 44492
rect 11655 44489 11667 44523
rect 11609 44483 11667 44489
rect 2608 44424 4384 44452
rect 2317 44387 2375 44393
rect 2317 44353 2329 44387
rect 2363 44353 2375 44387
rect 2317 44347 2375 44353
rect 2608 44316 2636 44424
rect 3050 44384 3056 44396
rect 3011 44356 3056 44384
rect 3050 44344 3056 44356
rect 3108 44344 3114 44396
rect 3234 44384 3240 44396
rect 3195 44356 3240 44384
rect 3234 44344 3240 44356
rect 3292 44344 3298 44396
rect 3697 44387 3755 44393
rect 3697 44353 3709 44387
rect 3743 44353 3755 44387
rect 3697 44347 3755 44353
rect 2240 44288 2636 44316
rect 3068 44316 3096 44344
rect 3326 44316 3332 44328
rect 3068 44288 3332 44316
rect 3326 44276 3332 44288
rect 3384 44316 3390 44328
rect 3712 44316 3740 44347
rect 3786 44344 3792 44396
rect 3844 44384 3850 44396
rect 4356 44393 4384 44424
rect 3881 44387 3939 44393
rect 3881 44384 3893 44387
rect 3844 44356 3893 44384
rect 3844 44344 3850 44356
rect 3881 44353 3893 44356
rect 3927 44353 3939 44387
rect 3881 44347 3939 44353
rect 4341 44387 4399 44393
rect 4341 44353 4353 44387
rect 4387 44353 4399 44387
rect 4341 44347 4399 44353
rect 3384 44288 3740 44316
rect 3896 44316 3924 44347
rect 4430 44344 4436 44396
rect 4488 44384 4494 44396
rect 4525 44387 4583 44393
rect 4525 44384 4537 44387
rect 4488 44356 4537 44384
rect 4488 44344 4494 44356
rect 4525 44353 4537 44356
rect 4571 44353 4583 44387
rect 4525 44347 4583 44353
rect 5258 44316 5264 44328
rect 3896 44288 5264 44316
rect 3384 44276 3390 44288
rect 5258 44276 5264 44288
rect 5316 44276 5322 44328
rect 983 44220 1716 44248
rect 1765 44251 1823 44257
rect 983 44217 995 44220
rect 937 44211 995 44217
rect 1765 44217 1777 44251
rect 1811 44248 1823 44251
rect 1811 44220 2774 44248
rect 1811 44217 1823 44220
rect 1765 44211 1823 44217
rect 658 44140 664 44192
rect 716 44180 722 44192
rect 1118 44180 1124 44192
rect 716 44152 1124 44180
rect 716 44140 722 44152
rect 1118 44140 1124 44152
rect 1176 44140 1182 44192
rect 2406 44140 2412 44192
rect 2464 44180 2470 44192
rect 2501 44183 2559 44189
rect 2501 44180 2513 44183
rect 2464 44152 2513 44180
rect 2464 44140 2470 44152
rect 2501 44149 2513 44152
rect 2547 44149 2559 44183
rect 2746 44180 2774 44220
rect 3878 44208 3884 44260
rect 3936 44248 3942 44260
rect 4430 44248 4436 44260
rect 3936 44220 4436 44248
rect 3936 44208 3942 44220
rect 4430 44208 4436 44220
rect 4488 44208 4494 44260
rect 5442 44180 5448 44192
rect 2746 44152 5448 44180
rect 2501 44143 2559 44149
rect 5442 44140 5448 44152
rect 5500 44140 5506 44192
rect 1104 44090 10856 44112
rect 106 44004 112 44056
rect 164 44044 170 44056
rect 658 44044 664 44056
rect 164 44016 664 44044
rect 164 44004 170 44016
rect 658 44004 664 44016
rect 716 44004 722 44056
rect 1104 44038 2582 44090
rect 2634 44038 2646 44090
rect 2698 44038 2710 44090
rect 2762 44038 2774 44090
rect 2826 44038 2838 44090
rect 2890 44038 5845 44090
rect 5897 44038 5909 44090
rect 5961 44038 5973 44090
rect 6025 44038 6037 44090
rect 6089 44038 6101 44090
rect 6153 44038 9109 44090
rect 9161 44038 9173 44090
rect 9225 44038 9237 44090
rect 9289 44038 9301 44090
rect 9353 44038 9365 44090
rect 9417 44038 10856 44090
rect 1104 44016 10856 44038
rect 1578 43976 1584 43988
rect 1539 43948 1584 43976
rect 1578 43936 1584 43948
rect 1636 43936 1642 43988
rect 8294 43976 8300 43988
rect 2746 43948 8300 43976
rect 1394 43772 1400 43784
rect 1355 43744 1400 43772
rect 1394 43732 1400 43744
rect 1452 43732 1458 43784
rect 2222 43732 2228 43784
rect 2280 43732 2286 43784
rect 2409 43775 2467 43781
rect 2409 43741 2421 43775
rect 2455 43772 2467 43775
rect 2746 43772 2774 43948
rect 8294 43936 8300 43948
rect 8352 43936 8358 43988
rect 4430 43908 4436 43920
rect 4391 43880 4436 43908
rect 4430 43868 4436 43880
rect 4488 43868 4494 43920
rect 3602 43840 3608 43852
rect 2884 43812 3608 43840
rect 2884 43781 2912 43812
rect 3602 43800 3608 43812
rect 3660 43800 3666 43852
rect 2455 43744 2774 43772
rect 2869 43775 2927 43781
rect 2455 43741 2467 43744
rect 2409 43735 2467 43741
rect 2869 43741 2881 43775
rect 2915 43741 2927 43775
rect 2869 43735 2927 43741
rect 3418 43732 3424 43784
rect 3476 43772 3482 43784
rect 4249 43775 4307 43781
rect 4249 43772 4261 43775
rect 3476 43744 4261 43772
rect 3476 43732 3482 43744
rect 4249 43741 4261 43744
rect 4295 43741 4307 43775
rect 4249 43735 4307 43741
rect 4893 43775 4951 43781
rect 4893 43741 4905 43775
rect 4939 43741 4951 43775
rect 5074 43772 5080 43784
rect 5035 43744 5080 43772
rect 4893 43735 4951 43741
rect 1762 43664 1768 43716
rect 1820 43704 1826 43716
rect 2240 43704 2268 43732
rect 1820 43676 2268 43704
rect 4908 43704 4936 43735
rect 5074 43732 5080 43744
rect 5132 43732 5138 43784
rect 9858 43772 9864 43784
rect 9819 43744 9864 43772
rect 9858 43732 9864 43744
rect 9916 43732 9922 43784
rect 5442 43704 5448 43716
rect 4908 43676 5448 43704
rect 1820 43664 1826 43676
rect 5442 43664 5448 43676
rect 5500 43664 5506 43716
rect 2222 43636 2228 43648
rect 2183 43608 2228 43636
rect 2222 43596 2228 43608
rect 2280 43596 2286 43648
rect 3050 43636 3056 43648
rect 3011 43608 3056 43636
rect 3050 43596 3056 43608
rect 3108 43596 3114 43648
rect 4985 43639 5043 43645
rect 4985 43605 4997 43639
rect 5031 43636 5043 43639
rect 9858 43636 9864 43648
rect 5031 43608 9864 43636
rect 5031 43605 5043 43608
rect 4985 43599 5043 43605
rect 9858 43596 9864 43608
rect 9916 43596 9922 43648
rect 10042 43636 10048 43648
rect 10003 43608 10048 43636
rect 10042 43596 10048 43608
rect 10100 43596 10106 43648
rect 1104 43546 10856 43568
rect 1104 43494 4213 43546
rect 4265 43494 4277 43546
rect 4329 43494 4341 43546
rect 4393 43494 4405 43546
rect 4457 43494 4469 43546
rect 4521 43494 7477 43546
rect 7529 43494 7541 43546
rect 7593 43494 7605 43546
rect 7657 43494 7669 43546
rect 7721 43494 7733 43546
rect 7785 43494 10856 43546
rect 1104 43472 10856 43494
rect 934 43392 940 43444
rect 992 43432 998 43444
rect 2225 43435 2283 43441
rect 2225 43432 2237 43435
rect 992 43404 2237 43432
rect 992 43392 998 43404
rect 2225 43401 2237 43404
rect 2271 43401 2283 43435
rect 2225 43395 2283 43401
rect 2148 43336 2774 43364
rect 1673 43299 1731 43305
rect 1673 43265 1685 43299
rect 1719 43296 1731 43299
rect 1762 43296 1768 43308
rect 1719 43268 1768 43296
rect 1719 43265 1731 43268
rect 1673 43259 1731 43265
rect 1762 43256 1768 43268
rect 1820 43256 1826 43308
rect 2148 43305 2176 43336
rect 2133 43299 2191 43305
rect 2133 43265 2145 43299
rect 2179 43265 2191 43299
rect 2133 43259 2191 43265
rect 2317 43299 2375 43305
rect 2317 43265 2329 43299
rect 2363 43265 2375 43299
rect 2746 43296 2774 43336
rect 3053 43299 3111 43305
rect 3053 43296 3065 43299
rect 2746 43268 3065 43296
rect 2317 43259 2375 43265
rect 3053 43265 3065 43268
rect 3099 43296 3111 43299
rect 3326 43296 3332 43308
rect 3099 43268 3332 43296
rect 3099 43265 3111 43268
rect 3053 43259 3111 43265
rect 1486 43188 1492 43240
rect 1544 43188 1550 43240
rect 1504 43160 1532 43188
rect 1762 43160 1768 43172
rect 1504 43132 1768 43160
rect 1762 43120 1768 43132
rect 1820 43120 1826 43172
rect 1486 43092 1492 43104
rect 1447 43064 1492 43092
rect 1486 43052 1492 43064
rect 1544 43052 1550 43104
rect 2332 43092 2360 43259
rect 3326 43256 3332 43268
rect 3384 43256 3390 43308
rect 9858 43296 9864 43308
rect 9819 43268 9864 43296
rect 9858 43256 9864 43268
rect 9916 43256 9922 43308
rect 2777 43231 2835 43237
rect 2777 43197 2789 43231
rect 2823 43228 2835 43231
rect 2866 43228 2872 43240
rect 2823 43200 2872 43228
rect 2823 43197 2835 43200
rect 2777 43191 2835 43197
rect 2866 43188 2872 43200
rect 2924 43188 2930 43240
rect 5442 43092 5448 43104
rect 2332 43064 5448 43092
rect 5442 43052 5448 43064
rect 5500 43052 5506 43104
rect 10042 43092 10048 43104
rect 10003 43064 10048 43092
rect 10042 43052 10048 43064
rect 10100 43052 10106 43104
rect 1104 43002 10856 43024
rect 1104 42950 2582 43002
rect 2634 42950 2646 43002
rect 2698 42950 2710 43002
rect 2762 42950 2774 43002
rect 2826 42950 2838 43002
rect 2890 42950 5845 43002
rect 5897 42950 5909 43002
rect 5961 42950 5973 43002
rect 6025 42950 6037 43002
rect 6089 42950 6101 43002
rect 6153 42950 9109 43002
rect 9161 42950 9173 43002
rect 9225 42950 9237 43002
rect 9289 42950 9301 43002
rect 9353 42950 9365 43002
rect 9417 42950 10856 43002
rect 1104 42928 10856 42950
rect 2130 42848 2136 42900
rect 2188 42888 2194 42900
rect 3326 42888 3332 42900
rect 2188 42860 3332 42888
rect 2188 42848 2194 42860
rect 3326 42848 3332 42860
rect 3384 42848 3390 42900
rect 4522 42820 4528 42832
rect 1688 42792 4528 42820
rect 1688 42693 1716 42792
rect 4522 42780 4528 42792
rect 4580 42780 4586 42832
rect 1673 42687 1731 42693
rect 1673 42653 1685 42687
rect 1719 42653 1731 42687
rect 1673 42647 1731 42653
rect 2314 42644 2320 42696
rect 2372 42684 2378 42696
rect 2409 42687 2467 42693
rect 2409 42684 2421 42687
rect 2372 42656 2421 42684
rect 2372 42644 2378 42656
rect 2409 42653 2421 42656
rect 2455 42653 2467 42687
rect 9858 42684 9864 42696
rect 9819 42656 9864 42684
rect 2409 42647 2467 42653
rect 9858 42644 9864 42656
rect 9916 42644 9922 42696
rect 1394 42508 1400 42560
rect 1452 42548 1458 42560
rect 1489 42551 1547 42557
rect 1489 42548 1501 42551
rect 1452 42520 1501 42548
rect 1452 42508 1458 42520
rect 1489 42517 1501 42520
rect 1535 42517 1547 42551
rect 2222 42548 2228 42560
rect 2183 42520 2228 42548
rect 1489 42511 1547 42517
rect 2222 42508 2228 42520
rect 2280 42508 2286 42560
rect 10042 42548 10048 42560
rect 10003 42520 10048 42548
rect 10042 42508 10048 42520
rect 10100 42508 10106 42560
rect 1104 42458 10856 42480
rect 1104 42406 4213 42458
rect 4265 42406 4277 42458
rect 4329 42406 4341 42458
rect 4393 42406 4405 42458
rect 4457 42406 4469 42458
rect 4521 42406 7477 42458
rect 7529 42406 7541 42458
rect 7593 42406 7605 42458
rect 7657 42406 7669 42458
rect 7721 42406 7733 42458
rect 7785 42406 10856 42458
rect 1104 42384 10856 42406
rect 5718 42344 5724 42356
rect 1688 42316 5724 42344
rect 1688 42217 1716 42316
rect 5718 42304 5724 42316
rect 5776 42304 5782 42356
rect 3418 42276 3424 42288
rect 3379 42248 3424 42276
rect 3418 42236 3424 42248
rect 3476 42276 3482 42288
rect 3602 42276 3608 42288
rect 3476 42248 3608 42276
rect 3476 42236 3482 42248
rect 3602 42236 3608 42248
rect 3660 42276 3666 42288
rect 4157 42279 4215 42285
rect 4157 42276 4169 42279
rect 3660 42248 4169 42276
rect 3660 42236 3666 42248
rect 4157 42245 4169 42248
rect 4203 42245 4215 42279
rect 4338 42276 4344 42288
rect 4251 42248 4344 42276
rect 4157 42239 4215 42245
rect 4338 42236 4344 42248
rect 4396 42276 4402 42288
rect 5074 42276 5080 42288
rect 4396 42248 5080 42276
rect 4396 42236 4402 42248
rect 5074 42236 5080 42248
rect 5132 42236 5138 42288
rect 1673 42211 1731 42217
rect 1673 42177 1685 42211
rect 1719 42177 1731 42211
rect 1673 42171 1731 42177
rect 4522 42168 4528 42220
rect 4580 42208 4586 42220
rect 4982 42208 4988 42220
rect 4580 42180 4988 42208
rect 4580 42168 4586 42180
rect 4982 42168 4988 42180
rect 5040 42168 5046 42220
rect 3605 42075 3663 42081
rect 3605 42041 3617 42075
rect 3651 42072 3663 42075
rect 3970 42072 3976 42084
rect 3651 42044 3976 42072
rect 3651 42041 3663 42044
rect 3605 42035 3663 42041
rect 3970 42032 3976 42044
rect 4028 42032 4034 42084
rect 1486 42004 1492 42016
rect 1447 41976 1492 42004
rect 1486 41964 1492 41976
rect 1544 41964 1550 42016
rect 1104 41914 10856 41936
rect 1104 41862 2582 41914
rect 2634 41862 2646 41914
rect 2698 41862 2710 41914
rect 2762 41862 2774 41914
rect 2826 41862 2838 41914
rect 2890 41862 5845 41914
rect 5897 41862 5909 41914
rect 5961 41862 5973 41914
rect 6025 41862 6037 41914
rect 6089 41862 6101 41914
rect 6153 41862 9109 41914
rect 9161 41862 9173 41914
rect 9225 41862 9237 41914
rect 9289 41862 9301 41914
rect 9353 41862 9365 41914
rect 9417 41862 10856 41914
rect 1104 41840 10856 41862
rect 1302 41760 1308 41812
rect 1360 41800 1366 41812
rect 2133 41803 2191 41809
rect 2133 41800 2145 41803
rect 1360 41772 2145 41800
rect 1360 41760 1366 41772
rect 2133 41769 2145 41772
rect 2179 41769 2191 41803
rect 2133 41763 2191 41769
rect 4065 41803 4123 41809
rect 4065 41769 4077 41803
rect 4111 41800 4123 41803
rect 9858 41800 9864 41812
rect 4111 41772 9864 41800
rect 4111 41769 4123 41772
rect 4065 41763 4123 41769
rect 9858 41760 9864 41772
rect 9916 41760 9922 41812
rect 4154 41664 4160 41676
rect 1688 41636 4160 41664
rect 1688 41605 1716 41636
rect 4154 41624 4160 41636
rect 4212 41624 4218 41676
rect 4614 41624 4620 41676
rect 4672 41664 4678 41676
rect 4672 41636 4844 41664
rect 4672 41624 4678 41636
rect 4816 41608 4844 41636
rect 1673 41599 1731 41605
rect 1673 41565 1685 41599
rect 1719 41565 1731 41599
rect 1673 41559 1731 41565
rect 1762 41556 1768 41608
rect 1820 41596 1826 41608
rect 2317 41599 2375 41605
rect 2317 41596 2329 41599
rect 1820 41568 2329 41596
rect 1820 41556 1826 41568
rect 2317 41565 2329 41568
rect 2363 41565 2375 41599
rect 3234 41596 3240 41608
rect 2317 41559 2375 41565
rect 2746 41568 3240 41596
rect 1026 41488 1032 41540
rect 1084 41528 1090 41540
rect 2746 41528 2774 41568
rect 3234 41556 3240 41568
rect 3292 41596 3298 41608
rect 3881 41599 3939 41605
rect 3881 41596 3893 41599
rect 3292 41568 3893 41596
rect 3292 41556 3298 41568
rect 3881 41565 3893 41568
rect 3927 41565 3939 41599
rect 3881 41559 3939 41565
rect 4065 41599 4123 41605
rect 4065 41565 4077 41599
rect 4111 41596 4123 41599
rect 4338 41596 4344 41608
rect 4111 41568 4344 41596
rect 4111 41565 4123 41568
rect 4065 41559 4123 41565
rect 4338 41556 4344 41568
rect 4396 41556 4402 41608
rect 4798 41556 4804 41608
rect 4856 41556 4862 41608
rect 5626 41556 5632 41608
rect 5684 41596 5690 41608
rect 6362 41596 6368 41608
rect 5684 41568 6368 41596
rect 5684 41556 5690 41568
rect 6362 41556 6368 41568
rect 6420 41556 6426 41608
rect 9861 41599 9919 41605
rect 9861 41565 9873 41599
rect 9907 41596 9919 41599
rect 11057 41599 11115 41605
rect 11057 41596 11069 41599
rect 9907 41568 11069 41596
rect 9907 41565 9919 41568
rect 9861 41559 9919 41565
rect 11057 41565 11069 41568
rect 11103 41565 11115 41599
rect 11057 41559 11115 41565
rect 6454 41528 6460 41540
rect 1084 41500 2774 41528
rect 5736 41500 6460 41528
rect 1084 41488 1090 41500
rect 5736 41472 5764 41500
rect 6454 41488 6460 41500
rect 6512 41488 6518 41540
rect 1394 41420 1400 41472
rect 1452 41460 1458 41472
rect 1489 41463 1547 41469
rect 1489 41460 1501 41463
rect 1452 41432 1501 41460
rect 1452 41420 1458 41432
rect 1489 41429 1501 41432
rect 1535 41429 1547 41463
rect 1489 41423 1547 41429
rect 3694 41420 3700 41472
rect 3752 41460 3758 41472
rect 5350 41460 5356 41472
rect 3752 41432 5356 41460
rect 3752 41420 3758 41432
rect 5350 41420 5356 41432
rect 5408 41420 5414 41472
rect 5718 41420 5724 41472
rect 5776 41420 5782 41472
rect 6086 41420 6092 41472
rect 6144 41460 6150 41472
rect 6362 41460 6368 41472
rect 6144 41432 6368 41460
rect 6144 41420 6150 41432
rect 6362 41420 6368 41432
rect 6420 41420 6426 41472
rect 10042 41460 10048 41472
rect 10003 41432 10048 41460
rect 10042 41420 10048 41432
rect 10100 41420 10106 41472
rect 1104 41370 10856 41392
rect 1104 41318 4213 41370
rect 4265 41318 4277 41370
rect 4329 41318 4341 41370
rect 4393 41318 4405 41370
rect 4457 41318 4469 41370
rect 4521 41318 7477 41370
rect 7529 41318 7541 41370
rect 7593 41318 7605 41370
rect 7657 41318 7669 41370
rect 7721 41318 7733 41370
rect 7785 41318 10856 41370
rect 1104 41296 10856 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 1670 41256 1676 41268
rect 1636 41228 1676 41256
rect 1636 41216 1642 41228
rect 1670 41216 1676 41228
rect 1728 41216 1734 41268
rect 1765 41259 1823 41265
rect 1765 41225 1777 41259
rect 1811 41256 1823 41259
rect 6270 41256 6276 41268
rect 1811 41228 6276 41256
rect 1811 41225 1823 41228
rect 1765 41219 1823 41225
rect 6270 41216 6276 41228
rect 6328 41216 6334 41268
rect 937 41191 995 41197
rect 937 41157 949 41191
rect 983 41188 995 41191
rect 983 41160 1808 41188
rect 983 41157 995 41160
rect 937 41151 995 41157
rect 1780 41132 1808 41160
rect 2222 41148 2228 41200
rect 2280 41148 2286 41200
rect 11885 41191 11943 41197
rect 11885 41188 11897 41191
rect 2746 41160 11897 41188
rect 1486 41120 1492 41132
rect 1447 41092 1492 41120
rect 1486 41080 1492 41092
rect 1544 41080 1550 41132
rect 1762 41120 1768 41132
rect 1723 41092 1768 41120
rect 1762 41080 1768 41092
rect 1820 41080 1826 41132
rect 1504 41052 1532 41080
rect 2240 41052 2268 41148
rect 2593 41123 2651 41129
rect 2593 41089 2605 41123
rect 2639 41120 2651 41123
rect 2746 41120 2774 41160
rect 11885 41157 11897 41160
rect 11931 41157 11943 41191
rect 11885 41151 11943 41157
rect 2639 41092 2774 41120
rect 2639 41089 2651 41092
rect 2593 41083 2651 41089
rect 5534 41080 5540 41132
rect 5592 41120 5598 41132
rect 6270 41120 6276 41132
rect 5592 41092 6276 41120
rect 5592 41080 5598 41092
rect 6270 41080 6276 41092
rect 6328 41080 6334 41132
rect 9858 41120 9864 41132
rect 9819 41092 9864 41120
rect 9858 41080 9864 41092
rect 9916 41080 9922 41132
rect 1504 41024 2268 41052
rect 2314 40944 2320 40996
rect 2372 40984 2378 40996
rect 2409 40987 2467 40993
rect 2409 40984 2421 40987
rect 2372 40956 2421 40984
rect 2372 40944 2378 40956
rect 2409 40953 2421 40956
rect 2455 40953 2467 40987
rect 2409 40947 2467 40953
rect 5534 40944 5540 40996
rect 5592 40984 5598 40996
rect 5902 40984 5908 40996
rect 5592 40956 5908 40984
rect 5592 40944 5598 40956
rect 5902 40944 5908 40956
rect 5960 40944 5966 40996
rect 10042 40916 10048 40928
rect 10003 40888 10048 40916
rect 10042 40876 10048 40888
rect 10100 40876 10106 40928
rect 1104 40826 10856 40848
rect 1104 40774 2582 40826
rect 2634 40774 2646 40826
rect 2698 40774 2710 40826
rect 2762 40774 2774 40826
rect 2826 40774 2838 40826
rect 2890 40774 5845 40826
rect 5897 40774 5909 40826
rect 5961 40774 5973 40826
rect 6025 40774 6037 40826
rect 6089 40774 6101 40826
rect 6153 40774 9109 40826
rect 9161 40774 9173 40826
rect 9225 40774 9237 40826
rect 9289 40774 9301 40826
rect 9353 40774 9365 40826
rect 9417 40774 10856 40826
rect 1104 40752 10856 40774
rect 3786 40712 3792 40724
rect 3747 40684 3792 40712
rect 3786 40672 3792 40684
rect 3844 40672 3850 40724
rect 3326 40604 3332 40656
rect 3384 40644 3390 40656
rect 3510 40644 3516 40656
rect 3384 40616 3516 40644
rect 3384 40604 3390 40616
rect 3510 40604 3516 40616
rect 3568 40604 3574 40656
rect 2774 40536 2780 40588
rect 2832 40576 2838 40588
rect 3050 40576 3056 40588
rect 2832 40548 3056 40576
rect 2832 40536 2838 40548
rect 3050 40536 3056 40548
rect 3108 40536 3114 40588
rect 11149 40579 11207 40585
rect 11149 40576 11161 40579
rect 3436 40548 11161 40576
rect 1670 40508 1676 40520
rect 1631 40480 1676 40508
rect 1670 40468 1676 40480
rect 1728 40468 1734 40520
rect 2133 40511 2191 40517
rect 2133 40477 2145 40511
rect 2179 40508 2191 40511
rect 2869 40511 2927 40517
rect 2179 40480 2774 40508
rect 2179 40477 2191 40480
rect 2133 40471 2191 40477
rect 2746 40440 2774 40480
rect 2869 40477 2881 40511
rect 2915 40508 2927 40511
rect 3436 40508 3464 40548
rect 11149 40545 11161 40548
rect 11195 40545 11207 40579
rect 11149 40539 11207 40545
rect 2915 40480 3464 40508
rect 2915 40477 2927 40480
rect 2869 40471 2927 40477
rect 3510 40468 3516 40520
rect 3568 40508 3574 40520
rect 3789 40511 3847 40517
rect 3789 40508 3801 40511
rect 3568 40480 3801 40508
rect 3568 40468 3574 40480
rect 3789 40477 3801 40480
rect 3835 40477 3847 40511
rect 3789 40471 3847 40477
rect 3973 40511 4031 40517
rect 3973 40477 3985 40511
rect 4019 40477 4031 40511
rect 3973 40471 4031 40477
rect 2746 40412 3188 40440
rect 1486 40372 1492 40384
rect 1447 40344 1492 40372
rect 1486 40332 1492 40344
rect 1544 40332 1550 40384
rect 1670 40332 1676 40384
rect 1728 40372 1734 40384
rect 1854 40372 1860 40384
rect 1728 40344 1860 40372
rect 1728 40332 1734 40344
rect 1854 40332 1860 40344
rect 1912 40332 1918 40384
rect 2314 40372 2320 40384
rect 2275 40344 2320 40372
rect 2314 40332 2320 40344
rect 2372 40332 2378 40384
rect 3050 40372 3056 40384
rect 3011 40344 3056 40372
rect 3050 40332 3056 40344
rect 3108 40332 3114 40384
rect 3160 40372 3188 40412
rect 3694 40400 3700 40452
rect 3752 40440 3758 40452
rect 3988 40440 4016 40471
rect 3752 40412 4016 40440
rect 3752 40400 3758 40412
rect 11701 40375 11759 40381
rect 11701 40372 11713 40375
rect 3160 40344 11713 40372
rect 11701 40341 11713 40344
rect 11747 40341 11759 40375
rect 11701 40335 11759 40341
rect 1104 40282 10856 40304
rect 1104 40230 4213 40282
rect 4265 40230 4277 40282
rect 4329 40230 4341 40282
rect 4393 40230 4405 40282
rect 4457 40230 4469 40282
rect 4521 40230 7477 40282
rect 7529 40230 7541 40282
rect 7593 40230 7605 40282
rect 7657 40230 7669 40282
rect 7721 40230 7733 40282
rect 7785 40230 10856 40282
rect 1104 40208 10856 40230
rect 750 40128 756 40180
rect 808 40168 814 40180
rect 1949 40171 2007 40177
rect 1949 40168 1961 40171
rect 808 40140 1961 40168
rect 808 40128 814 40140
rect 1949 40137 1961 40140
rect 1995 40137 2007 40171
rect 1949 40131 2007 40137
rect 2774 40100 2780 40112
rect 2735 40072 2780 40100
rect 2774 40060 2780 40072
rect 2832 40100 2838 40112
rect 3234 40100 3240 40112
rect 2832 40072 3240 40100
rect 2832 40060 2838 40072
rect 3234 40060 3240 40072
rect 3292 40060 3298 40112
rect 3970 40060 3976 40112
rect 4028 40100 4034 40112
rect 4028 40072 4292 40100
rect 4028 40060 4034 40072
rect 1854 39992 1860 40044
rect 1912 40032 1918 40044
rect 1949 40035 2007 40041
rect 1949 40032 1961 40035
rect 1912 40004 1961 40032
rect 1912 39992 1918 40004
rect 1949 40001 1961 40004
rect 1995 40001 2007 40035
rect 1949 39995 2007 40001
rect 2225 40035 2283 40041
rect 2225 40001 2237 40035
rect 2271 40032 2283 40035
rect 2866 40032 2872 40044
rect 2271 40004 2872 40032
rect 2271 40001 2283 40004
rect 2225 39995 2283 40001
rect 1964 39964 1992 39995
rect 2866 39992 2872 40004
rect 2924 39992 2930 40044
rect 2961 40035 3019 40041
rect 2961 40001 2973 40035
rect 3007 40032 3019 40035
rect 3421 40035 3479 40041
rect 3421 40032 3433 40035
rect 3007 40004 3433 40032
rect 3007 40001 3019 40004
rect 2961 39995 3019 40001
rect 3421 40001 3433 40004
rect 3467 40032 3479 40035
rect 3510 40032 3516 40044
rect 3467 40004 3516 40032
rect 3467 40001 3479 40004
rect 3421 39995 3479 40001
rect 2976 39964 3004 39995
rect 3510 39992 3516 40004
rect 3568 39992 3574 40044
rect 3605 40035 3663 40041
rect 3605 40001 3617 40035
rect 3651 40032 3663 40035
rect 3786 40032 3792 40044
rect 3651 40004 3792 40032
rect 3651 40001 3663 40004
rect 3605 39995 3663 40001
rect 3786 39992 3792 40004
rect 3844 40032 3850 40044
rect 4264 40041 4292 40072
rect 4071 40035 4129 40041
rect 4071 40032 4083 40035
rect 3844 40004 4083 40032
rect 3844 39992 3850 40004
rect 4071 40001 4083 40004
rect 4117 40001 4129 40035
rect 4071 39995 4129 40001
rect 4249 40035 4307 40041
rect 4249 40001 4261 40035
rect 4295 40032 4307 40035
rect 4522 40032 4528 40044
rect 4295 40004 4528 40032
rect 4295 40001 4307 40004
rect 4249 39995 4307 40001
rect 4522 39992 4528 40004
rect 4580 39992 4586 40044
rect 9861 40035 9919 40041
rect 9861 40001 9873 40035
rect 9907 40001 9919 40035
rect 9861 39995 9919 40001
rect 1964 39936 3004 39964
rect 4157 39967 4215 39973
rect 4157 39933 4169 39967
rect 4203 39964 4215 39967
rect 9876 39964 9904 39995
rect 4203 39936 9904 39964
rect 4203 39933 4215 39936
rect 4157 39927 4215 39933
rect 2866 39856 2872 39908
rect 2924 39856 2930 39908
rect 3421 39899 3479 39905
rect 3421 39865 3433 39899
rect 3467 39896 3479 39899
rect 5166 39896 5172 39908
rect 3467 39868 5172 39896
rect 3467 39865 3479 39868
rect 3421 39859 3479 39865
rect 5166 39856 5172 39868
rect 5224 39856 5230 39908
rect 10042 39896 10048 39908
rect 10003 39868 10048 39896
rect 10042 39856 10048 39868
rect 10100 39856 10106 39908
rect 2884 39828 2912 39856
rect 3878 39828 3884 39840
rect 2884 39800 3884 39828
rect 3878 39788 3884 39800
rect 3936 39788 3942 39840
rect 4338 39788 4344 39840
rect 4396 39828 4402 39840
rect 8478 39828 8484 39840
rect 4396 39800 8484 39828
rect 4396 39788 4402 39800
rect 8478 39788 8484 39800
rect 8536 39788 8542 39840
rect 1104 39738 10856 39760
rect 1104 39686 2582 39738
rect 2634 39686 2646 39738
rect 2698 39686 2710 39738
rect 2762 39686 2774 39738
rect 2826 39686 2838 39738
rect 2890 39686 5845 39738
rect 5897 39686 5909 39738
rect 5961 39686 5973 39738
rect 6025 39686 6037 39738
rect 6089 39686 6101 39738
rect 6153 39686 9109 39738
rect 9161 39686 9173 39738
rect 9225 39686 9237 39738
rect 9289 39686 9301 39738
rect 9353 39686 9365 39738
rect 9417 39686 10856 39738
rect 1104 39664 10856 39686
rect 3789 39627 3847 39633
rect 3789 39593 3801 39627
rect 3835 39624 3847 39627
rect 4890 39624 4896 39636
rect 3835 39596 4896 39624
rect 3835 39593 3847 39596
rect 3789 39587 3847 39593
rect 4890 39584 4896 39596
rect 4948 39584 4954 39636
rect 5166 39556 5172 39568
rect 2746 39528 5172 39556
rect 2746 39488 2774 39528
rect 5166 39516 5172 39528
rect 5224 39516 5230 39568
rect 4338 39488 4344 39500
rect 1688 39460 2774 39488
rect 3160 39460 4344 39488
rect 1688 39429 1716 39460
rect 1673 39423 1731 39429
rect 1673 39389 1685 39423
rect 1719 39389 1731 39423
rect 2406 39420 2412 39432
rect 2367 39392 2412 39420
rect 1673 39383 1731 39389
rect 2406 39380 2412 39392
rect 2464 39380 2470 39432
rect 3160 39429 3188 39460
rect 4338 39448 4344 39460
rect 4396 39448 4402 39500
rect 4525 39491 4583 39497
rect 4525 39457 4537 39491
rect 4571 39488 4583 39491
rect 4571 39460 9904 39488
rect 4571 39457 4583 39460
rect 4525 39451 4583 39457
rect 3145 39423 3203 39429
rect 3145 39389 3157 39423
rect 3191 39389 3203 39423
rect 3145 39383 3203 39389
rect 3789 39423 3847 39429
rect 3789 39389 3801 39423
rect 3835 39389 3847 39423
rect 3789 39383 3847 39389
rect 1854 39312 1860 39364
rect 1912 39352 1918 39364
rect 3804 39352 3832 39383
rect 3878 39380 3884 39432
rect 3936 39420 3942 39432
rect 3973 39423 4031 39429
rect 3973 39420 3985 39423
rect 3936 39392 3985 39420
rect 3936 39380 3942 39392
rect 3973 39389 3985 39392
rect 4019 39389 4031 39423
rect 3973 39383 4031 39389
rect 4062 39380 4068 39432
rect 4120 39420 4126 39432
rect 9876 39429 9904 39460
rect 4433 39423 4491 39429
rect 4433 39420 4445 39423
rect 4120 39392 4445 39420
rect 4120 39380 4126 39392
rect 4433 39389 4445 39392
rect 4479 39389 4491 39423
rect 4617 39423 4675 39429
rect 4617 39420 4629 39423
rect 4433 39383 4491 39389
rect 4540 39392 4629 39420
rect 4540 39364 4568 39392
rect 4617 39389 4629 39392
rect 4663 39389 4675 39423
rect 4617 39383 4675 39389
rect 9861 39423 9919 39429
rect 9861 39389 9873 39423
rect 9907 39389 9919 39423
rect 9861 39383 9919 39389
rect 1912 39324 3832 39352
rect 1912 39312 1918 39324
rect 4522 39312 4528 39364
rect 4580 39312 4586 39364
rect 1394 39244 1400 39296
rect 1452 39284 1458 39296
rect 1489 39287 1547 39293
rect 1489 39284 1501 39287
rect 1452 39256 1501 39284
rect 1452 39244 1458 39256
rect 1489 39253 1501 39256
rect 1535 39253 1547 39287
rect 2222 39284 2228 39296
rect 2183 39256 2228 39284
rect 1489 39247 1547 39253
rect 2222 39244 2228 39256
rect 2280 39244 2286 39296
rect 2958 39284 2964 39296
rect 2919 39256 2964 39284
rect 2958 39244 2964 39256
rect 3016 39244 3022 39296
rect 3786 39244 3792 39296
rect 3844 39284 3850 39296
rect 5166 39284 5172 39296
rect 3844 39256 5172 39284
rect 3844 39244 3850 39256
rect 5166 39244 5172 39256
rect 5224 39244 5230 39296
rect 10042 39284 10048 39296
rect 10003 39256 10048 39284
rect 10042 39244 10048 39256
rect 10100 39244 10106 39296
rect 1104 39194 10856 39216
rect 1104 39142 4213 39194
rect 4265 39142 4277 39194
rect 4329 39142 4341 39194
rect 4393 39142 4405 39194
rect 4457 39142 4469 39194
rect 4521 39142 7477 39194
rect 7529 39142 7541 39194
rect 7593 39142 7605 39194
rect 7657 39142 7669 39194
rect 7721 39142 7733 39194
rect 7785 39142 10856 39194
rect 1104 39120 10856 39142
rect 4062 39080 4068 39092
rect 3528 39052 4068 39080
rect 842 38972 848 39024
rect 900 39012 906 39024
rect 1673 39015 1731 39021
rect 1673 39012 1685 39015
rect 900 38984 1685 39012
rect 900 38972 906 38984
rect 1673 38981 1685 38984
rect 1719 38981 1731 39015
rect 1673 38975 1731 38981
rect 2406 38972 2412 39024
rect 2464 39012 2470 39024
rect 2464 38984 2774 39012
rect 2464 38972 2470 38984
rect 2746 38956 2774 38984
rect 1854 38944 1860 38956
rect 1815 38916 1860 38944
rect 1854 38904 1860 38916
rect 1912 38904 1918 38956
rect 2041 38947 2099 38953
rect 2041 38913 2053 38947
rect 2087 38913 2099 38947
rect 2746 38916 2780 38956
rect 2041 38907 2099 38913
rect 2056 38876 2084 38907
rect 2774 38904 2780 38916
rect 2832 38904 2838 38956
rect 2866 38904 2872 38956
rect 2924 38944 2930 38956
rect 2961 38947 3019 38953
rect 2961 38944 2973 38947
rect 2924 38916 2973 38944
rect 2924 38904 2930 38916
rect 2961 38913 2973 38916
rect 3007 38913 3019 38947
rect 2961 38907 3019 38913
rect 2406 38876 2412 38888
rect 2056 38848 2412 38876
rect 2406 38836 2412 38848
rect 2464 38876 2470 38888
rect 3528 38876 3556 39052
rect 4062 39040 4068 39052
rect 4120 39040 4126 39092
rect 4341 39083 4399 39089
rect 4341 39049 4353 39083
rect 4387 39080 4399 39083
rect 9858 39080 9864 39092
rect 4387 39052 9864 39080
rect 4387 39049 4399 39052
rect 4341 39043 4399 39049
rect 9858 39040 9864 39052
rect 9916 39040 9922 39092
rect 3694 38972 3700 39024
rect 3752 38972 3758 39024
rect 3605 38947 3663 38953
rect 3605 38913 3617 38947
rect 3651 38944 3663 38947
rect 3712 38944 3740 38972
rect 3651 38916 3740 38944
rect 3651 38913 3663 38916
rect 3605 38907 3663 38913
rect 3786 38904 3792 38956
rect 3844 38944 3850 38956
rect 3970 38944 3976 38956
rect 3844 38916 3976 38944
rect 3844 38904 3850 38916
rect 3970 38904 3976 38916
rect 4028 38904 4034 38956
rect 4062 38904 4068 38956
rect 4120 38944 4126 38956
rect 4249 38947 4307 38953
rect 4249 38944 4261 38947
rect 4120 38916 4261 38944
rect 4120 38904 4126 38916
rect 4249 38913 4261 38916
rect 4295 38913 4307 38947
rect 4249 38907 4307 38913
rect 4430 38904 4436 38956
rect 4488 38944 4494 38956
rect 4982 38944 4988 38956
rect 4488 38916 4988 38944
rect 4488 38904 4494 38916
rect 4982 38904 4988 38916
rect 5040 38904 5046 38956
rect 9861 38947 9919 38953
rect 9861 38913 9873 38947
rect 9907 38913 9919 38947
rect 9861 38907 9919 38913
rect 2464 38848 3556 38876
rect 3697 38879 3755 38885
rect 2464 38836 2470 38848
rect 3697 38845 3709 38879
rect 3743 38876 3755 38879
rect 9876 38876 9904 38907
rect 3743 38848 9904 38876
rect 3743 38845 3755 38848
rect 3697 38839 3755 38845
rect 845 38811 903 38817
rect 845 38777 857 38811
rect 891 38808 903 38811
rect 1854 38808 1860 38820
rect 891 38780 1860 38808
rect 891 38777 903 38780
rect 845 38771 903 38777
rect 1854 38768 1860 38780
rect 1912 38768 1918 38820
rect 2774 38768 2780 38820
rect 2832 38768 2838 38820
rect 3145 38811 3203 38817
rect 3145 38777 3157 38811
rect 3191 38808 3203 38811
rect 3602 38808 3608 38820
rect 3191 38780 3608 38808
rect 3191 38777 3203 38780
rect 3145 38771 3203 38777
rect 3602 38768 3608 38780
rect 3660 38768 3666 38820
rect 2792 38740 2820 38768
rect 7006 38740 7012 38752
rect 2792 38712 7012 38740
rect 7006 38700 7012 38712
rect 7064 38700 7070 38752
rect 10042 38740 10048 38752
rect 10003 38712 10048 38740
rect 10042 38700 10048 38712
rect 10100 38700 10106 38752
rect 1104 38650 10856 38672
rect 1104 38598 2582 38650
rect 2634 38598 2646 38650
rect 2698 38598 2710 38650
rect 2762 38598 2774 38650
rect 2826 38598 2838 38650
rect 2890 38598 5845 38650
rect 5897 38598 5909 38650
rect 5961 38598 5973 38650
rect 6025 38598 6037 38650
rect 6089 38598 6101 38650
rect 6153 38598 9109 38650
rect 9161 38598 9173 38650
rect 9225 38598 9237 38650
rect 9289 38598 9301 38650
rect 9353 38598 9365 38650
rect 9417 38598 10856 38650
rect 1104 38576 10856 38598
rect 2869 38539 2927 38545
rect 2869 38505 2881 38539
rect 2915 38536 2927 38539
rect 3234 38536 3240 38548
rect 2915 38508 3240 38536
rect 2915 38505 2927 38508
rect 2869 38499 2927 38505
rect 2225 38335 2283 38341
rect 2225 38301 2237 38335
rect 2271 38332 2283 38335
rect 2774 38332 2780 38344
rect 2271 38304 2780 38332
rect 2271 38301 2283 38304
rect 2225 38295 2283 38301
rect 2774 38292 2780 38304
rect 2832 38332 2838 38344
rect 2884 38332 2912 38499
rect 3234 38496 3240 38508
rect 3292 38496 3298 38548
rect 3973 38539 4031 38545
rect 3973 38505 3985 38539
rect 4019 38536 4031 38539
rect 11057 38539 11115 38545
rect 11057 38536 11069 38539
rect 4019 38508 11069 38536
rect 4019 38505 4031 38508
rect 3973 38499 4031 38505
rect 11057 38505 11069 38508
rect 11103 38505 11115 38539
rect 11057 38499 11115 38505
rect 3510 38468 3516 38480
rect 3252 38440 3516 38468
rect 3252 38412 3280 38440
rect 3510 38428 3516 38440
rect 3568 38428 3574 38480
rect 3234 38360 3240 38412
rect 3292 38360 3298 38412
rect 4338 38400 4344 38412
rect 3804 38372 4344 38400
rect 2832 38304 2925 38332
rect 2832 38292 2838 38304
rect 3510 38292 3516 38344
rect 3568 38332 3574 38344
rect 3804 38341 3832 38372
rect 4338 38360 4344 38372
rect 4396 38360 4402 38412
rect 3789 38335 3847 38341
rect 3789 38332 3801 38335
rect 3568 38304 3801 38332
rect 3568 38292 3574 38304
rect 3789 38301 3801 38304
rect 3835 38301 3847 38335
rect 3789 38295 3847 38301
rect 3973 38335 4031 38341
rect 3973 38301 3985 38335
rect 4019 38332 4031 38335
rect 4430 38332 4436 38344
rect 4019 38304 4436 38332
rect 4019 38301 4031 38304
rect 3973 38295 4031 38301
rect 4430 38292 4436 38304
rect 4488 38292 4494 38344
rect 2961 38267 3019 38273
rect 2961 38233 2973 38267
rect 3007 38264 3019 38267
rect 4982 38264 4988 38276
rect 3007 38236 4988 38264
rect 3007 38233 3019 38236
rect 2961 38227 3019 38233
rect 4982 38224 4988 38236
rect 5040 38224 5046 38276
rect 2130 38196 2136 38208
rect 2091 38168 2136 38196
rect 2130 38156 2136 38168
rect 2188 38156 2194 38208
rect 2222 38156 2228 38208
rect 2280 38196 2286 38208
rect 4062 38196 4068 38208
rect 2280 38168 4068 38196
rect 2280 38156 2286 38168
rect 4062 38156 4068 38168
rect 4120 38156 4126 38208
rect 1104 38106 10856 38128
rect 1104 38054 4213 38106
rect 4265 38054 4277 38106
rect 4329 38054 4341 38106
rect 4393 38054 4405 38106
rect 4457 38054 4469 38106
rect 4521 38054 7477 38106
rect 7529 38054 7541 38106
rect 7593 38054 7605 38106
rect 7657 38054 7669 38106
rect 7721 38054 7733 38106
rect 7785 38054 10856 38106
rect 1104 38032 10856 38054
rect 1762 37952 1768 38004
rect 1820 37992 1826 38004
rect 2317 37995 2375 38001
rect 2317 37992 2329 37995
rect 1820 37964 2329 37992
rect 1820 37952 1826 37964
rect 2317 37961 2329 37964
rect 2363 37961 2375 37995
rect 2317 37955 2375 37961
rect 5626 37924 5632 37936
rect 1688 37896 5632 37924
rect 1688 37865 1716 37896
rect 5626 37884 5632 37896
rect 5684 37884 5690 37936
rect 1673 37859 1731 37865
rect 1673 37825 1685 37859
rect 1719 37825 1731 37859
rect 1673 37819 1731 37825
rect 2501 37859 2559 37865
rect 2501 37825 2513 37859
rect 2547 37856 2559 37859
rect 2774 37856 2780 37868
rect 2547 37828 2780 37856
rect 2547 37825 2559 37828
rect 2501 37819 2559 37825
rect 2774 37816 2780 37828
rect 2832 37816 2838 37868
rect 9858 37856 9864 37868
rect 9819 37828 9864 37856
rect 9858 37816 9864 37828
rect 9916 37816 9922 37868
rect 2222 37680 2228 37732
rect 2280 37720 2286 37732
rect 7282 37720 7288 37732
rect 2280 37692 7288 37720
rect 2280 37680 2286 37692
rect 7282 37680 7288 37692
rect 7340 37680 7346 37732
rect 1486 37652 1492 37664
rect 1447 37624 1492 37652
rect 1486 37612 1492 37624
rect 1544 37612 1550 37664
rect 10042 37652 10048 37664
rect 10003 37624 10048 37652
rect 10042 37612 10048 37624
rect 10100 37612 10106 37664
rect 1104 37562 10856 37584
rect 1104 37510 2582 37562
rect 2634 37510 2646 37562
rect 2698 37510 2710 37562
rect 2762 37510 2774 37562
rect 2826 37510 2838 37562
rect 2890 37510 5845 37562
rect 5897 37510 5909 37562
rect 5961 37510 5973 37562
rect 6025 37510 6037 37562
rect 6089 37510 6101 37562
rect 6153 37510 9109 37562
rect 9161 37510 9173 37562
rect 9225 37510 9237 37562
rect 9289 37510 9301 37562
rect 9353 37510 9365 37562
rect 9417 37510 10856 37562
rect 1104 37488 10856 37510
rect 2314 37448 2320 37460
rect 2275 37420 2320 37448
rect 2314 37408 2320 37420
rect 2372 37408 2378 37460
rect 2130 37340 2136 37392
rect 2188 37340 2194 37392
rect 2148 37312 2176 37340
rect 2314 37312 2320 37324
rect 1688 37284 2320 37312
rect 1489 37247 1547 37253
rect 1489 37213 1501 37247
rect 1535 37244 1547 37247
rect 1578 37244 1584 37256
rect 1535 37216 1584 37244
rect 1535 37213 1547 37216
rect 1489 37207 1547 37213
rect 1578 37204 1584 37216
rect 1636 37204 1642 37256
rect 1688 37253 1716 37284
rect 2314 37272 2320 37284
rect 2372 37272 2378 37324
rect 2424 37284 2636 37312
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37213 1731 37247
rect 1673 37207 1731 37213
rect 2130 37204 2136 37256
rect 2188 37244 2194 37256
rect 2424 37244 2452 37284
rect 2188 37216 2452 37244
rect 2501 37247 2559 37253
rect 2188 37204 2194 37216
rect 2501 37213 2513 37247
rect 2547 37213 2559 37247
rect 2608 37244 2636 37284
rect 2961 37247 3019 37253
rect 2961 37244 2973 37247
rect 2608 37216 2973 37244
rect 2501 37207 2559 37213
rect 2961 37213 2973 37216
rect 3007 37213 3019 37247
rect 2961 37207 3019 37213
rect 3053 37247 3111 37253
rect 3053 37213 3065 37247
rect 3099 37244 3111 37247
rect 3418 37244 3424 37256
rect 3099 37216 3424 37244
rect 3099 37213 3111 37216
rect 3053 37207 3111 37213
rect 2516 37176 2544 37207
rect 3418 37204 3424 37216
rect 3476 37204 3482 37256
rect 3970 37204 3976 37256
rect 4028 37244 4034 37256
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 4028 37216 9873 37244
rect 4028 37204 4034 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 11333 37179 11391 37185
rect 11333 37176 11345 37179
rect 2516 37148 11345 37176
rect 11333 37145 11345 37148
rect 11379 37145 11391 37179
rect 11333 37139 11391 37145
rect 1670 37108 1676 37120
rect 1631 37080 1676 37108
rect 1670 37068 1676 37080
rect 1728 37068 1734 37120
rect 2774 37068 2780 37120
rect 2832 37108 2838 37120
rect 8754 37108 8760 37120
rect 2832 37080 8760 37108
rect 2832 37068 2838 37080
rect 8754 37068 8760 37080
rect 8812 37068 8818 37120
rect 10042 37108 10048 37120
rect 10003 37080 10048 37108
rect 10042 37068 10048 37080
rect 10100 37068 10106 37120
rect 1104 37018 10856 37040
rect 1104 36966 4213 37018
rect 4265 36966 4277 37018
rect 4329 36966 4341 37018
rect 4393 36966 4405 37018
rect 4457 36966 4469 37018
rect 4521 36966 7477 37018
rect 7529 36966 7541 37018
rect 7593 36966 7605 37018
rect 7657 36966 7669 37018
rect 7721 36966 7733 37018
rect 7785 36966 10856 37018
rect 1104 36944 10856 36966
rect 1670 36864 1676 36916
rect 1728 36904 1734 36916
rect 3697 36907 3755 36913
rect 1728 36876 3648 36904
rect 1728 36864 1734 36876
rect 3620 36836 3648 36876
rect 3697 36873 3709 36907
rect 3743 36904 3755 36907
rect 9858 36904 9864 36916
rect 3743 36876 9864 36904
rect 3743 36873 3755 36876
rect 3697 36867 3755 36873
rect 9858 36864 9864 36876
rect 9916 36864 9922 36916
rect 5534 36836 5540 36848
rect 3620 36808 5540 36836
rect 5534 36796 5540 36808
rect 5592 36796 5598 36848
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 2222 36768 2228 36780
rect 1719 36740 2228 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 2222 36728 2228 36740
rect 2280 36728 2286 36780
rect 2409 36771 2467 36777
rect 2409 36737 2421 36771
rect 2455 36768 2467 36771
rect 2774 36768 2780 36780
rect 2455 36740 2780 36768
rect 2455 36737 2467 36740
rect 2409 36731 2467 36737
rect 2774 36728 2780 36740
rect 2832 36728 2838 36780
rect 2869 36771 2927 36777
rect 2869 36737 2881 36771
rect 2915 36737 2927 36771
rect 2869 36731 2927 36737
rect 2884 36700 2912 36731
rect 3510 36728 3516 36780
rect 3568 36768 3574 36780
rect 3605 36771 3663 36777
rect 3605 36768 3617 36771
rect 3568 36740 3617 36768
rect 3568 36728 3574 36740
rect 3605 36737 3617 36740
rect 3651 36737 3663 36771
rect 3786 36768 3792 36780
rect 3747 36740 3792 36768
rect 3605 36731 3663 36737
rect 3786 36728 3792 36740
rect 3844 36728 3850 36780
rect 11241 36771 11299 36777
rect 11241 36768 11253 36771
rect 4632 36740 11253 36768
rect 2884 36672 3372 36700
rect 3050 36632 3056 36644
rect 3011 36604 3056 36632
rect 3050 36592 3056 36604
rect 3108 36592 3114 36644
rect 3344 36632 3372 36672
rect 4632 36632 4660 36740
rect 11241 36737 11253 36740
rect 11287 36737 11299 36771
rect 11241 36731 11299 36737
rect 4890 36660 4896 36712
rect 4948 36700 4954 36712
rect 5442 36700 5448 36712
rect 4948 36672 5448 36700
rect 4948 36660 4954 36672
rect 5442 36660 5448 36672
rect 5500 36660 5506 36712
rect 3344 36604 4660 36632
rect 198 36524 204 36576
rect 256 36564 262 36576
rect 934 36564 940 36576
rect 256 36536 940 36564
rect 256 36524 262 36536
rect 934 36524 940 36536
rect 992 36524 998 36576
rect 1394 36524 1400 36576
rect 1452 36564 1458 36576
rect 1489 36567 1547 36573
rect 1489 36564 1501 36567
rect 1452 36536 1501 36564
rect 1452 36524 1458 36536
rect 1489 36533 1501 36536
rect 1535 36533 1547 36567
rect 2222 36564 2228 36576
rect 2183 36536 2228 36564
rect 1489 36527 1547 36533
rect 2222 36524 2228 36536
rect 2280 36524 2286 36576
rect 5074 36524 5080 36576
rect 5132 36564 5138 36576
rect 5442 36564 5448 36576
rect 5132 36536 5448 36564
rect 5132 36524 5138 36536
rect 5442 36524 5448 36536
rect 5500 36524 5506 36576
rect 7926 36524 7932 36576
rect 7984 36564 7990 36576
rect 8110 36564 8116 36576
rect 7984 36536 8116 36564
rect 7984 36524 7990 36536
rect 8110 36524 8116 36536
rect 8168 36524 8174 36576
rect 1104 36474 10856 36496
rect 1104 36422 2582 36474
rect 2634 36422 2646 36474
rect 2698 36422 2710 36474
rect 2762 36422 2774 36474
rect 2826 36422 2838 36474
rect 2890 36422 5845 36474
rect 5897 36422 5909 36474
rect 5961 36422 5973 36474
rect 6025 36422 6037 36474
rect 6089 36422 6101 36474
rect 6153 36422 9109 36474
rect 9161 36422 9173 36474
rect 9225 36422 9237 36474
rect 9289 36422 9301 36474
rect 9353 36422 9365 36474
rect 9417 36422 10856 36474
rect 1104 36400 10856 36422
rect 3970 36360 3976 36372
rect 3931 36332 3976 36360
rect 3970 36320 3976 36332
rect 4028 36320 4034 36372
rect 5166 36320 5172 36372
rect 5224 36360 5230 36372
rect 5534 36360 5540 36372
rect 5224 36332 5540 36360
rect 5224 36320 5230 36332
rect 5534 36320 5540 36332
rect 5592 36320 5598 36372
rect 3418 36252 3424 36304
rect 3476 36292 3482 36304
rect 3786 36292 3792 36304
rect 3476 36264 3792 36292
rect 3476 36252 3482 36264
rect 3786 36252 3792 36264
rect 3844 36252 3850 36304
rect 8570 36224 8576 36236
rect 2746 36196 8576 36224
rect 1673 36159 1731 36165
rect 1673 36125 1685 36159
rect 1719 36156 1731 36159
rect 2746 36156 2774 36196
rect 8570 36184 8576 36196
rect 8628 36184 8634 36236
rect 1719 36128 2774 36156
rect 1719 36125 1731 36128
rect 1673 36119 1731 36125
rect 3510 36116 3516 36168
rect 3568 36156 3574 36168
rect 3789 36159 3847 36165
rect 3789 36156 3801 36159
rect 3568 36128 3801 36156
rect 3568 36116 3574 36128
rect 3789 36125 3801 36128
rect 3835 36125 3847 36159
rect 3789 36119 3847 36125
rect 3878 36116 3884 36168
rect 3936 36156 3942 36168
rect 3973 36159 4031 36165
rect 3973 36156 3985 36159
rect 3936 36128 3985 36156
rect 3936 36116 3942 36128
rect 3973 36125 3985 36128
rect 4019 36125 4031 36159
rect 9858 36156 9864 36168
rect 9819 36128 9864 36156
rect 3973 36119 4031 36125
rect 9858 36116 9864 36128
rect 9916 36116 9922 36168
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 10042 36020 10048 36032
rect 10003 35992 10048 36020
rect 10042 35980 10048 35992
rect 10100 35980 10106 36032
rect 1104 35930 10856 35952
rect 1104 35878 4213 35930
rect 4265 35878 4277 35930
rect 4329 35878 4341 35930
rect 4393 35878 4405 35930
rect 4457 35878 4469 35930
rect 4521 35878 7477 35930
rect 7529 35878 7541 35930
rect 7593 35878 7605 35930
rect 7657 35878 7669 35930
rect 7721 35878 7733 35930
rect 7785 35878 10856 35930
rect 1104 35856 10856 35878
rect 1765 35819 1823 35825
rect 1765 35785 1777 35819
rect 1811 35816 1823 35819
rect 6914 35816 6920 35828
rect 1811 35788 6920 35816
rect 1811 35785 1823 35788
rect 1765 35779 1823 35785
rect 6914 35776 6920 35788
rect 6972 35776 6978 35828
rect 2314 35748 2320 35760
rect 1596 35720 2320 35748
rect 1596 35689 1624 35720
rect 2314 35708 2320 35720
rect 2372 35708 2378 35760
rect 3510 35748 3516 35760
rect 2792 35720 3516 35748
rect 1581 35683 1639 35689
rect 1581 35649 1593 35683
rect 1627 35649 1639 35683
rect 1762 35680 1768 35692
rect 1723 35652 1768 35680
rect 1581 35643 1639 35649
rect 1762 35640 1768 35652
rect 1820 35640 1826 35692
rect 2406 35640 2412 35692
rect 2464 35680 2470 35692
rect 2792 35689 2820 35720
rect 3510 35708 3516 35720
rect 3568 35708 3574 35760
rect 2501 35683 2559 35689
rect 2501 35680 2513 35683
rect 2464 35652 2513 35680
rect 2464 35640 2470 35652
rect 2501 35649 2513 35652
rect 2547 35649 2559 35683
rect 2501 35643 2559 35649
rect 2777 35683 2835 35689
rect 2777 35649 2789 35683
rect 2823 35649 2835 35683
rect 2777 35643 2835 35649
rect 3421 35683 3479 35689
rect 3421 35649 3433 35683
rect 3467 35680 3479 35683
rect 3602 35680 3608 35692
rect 3467 35652 3608 35680
rect 3467 35649 3479 35652
rect 3421 35643 3479 35649
rect 3602 35640 3608 35652
rect 3660 35640 3666 35692
rect 9766 35640 9772 35692
rect 9824 35680 9830 35692
rect 9861 35683 9919 35689
rect 9861 35680 9873 35683
rect 9824 35652 9873 35680
rect 9824 35640 9830 35652
rect 9861 35649 9873 35652
rect 9907 35649 9919 35683
rect 9861 35643 9919 35649
rect 3697 35615 3755 35621
rect 3697 35581 3709 35615
rect 3743 35612 3755 35615
rect 4154 35612 4160 35624
rect 3743 35584 4160 35612
rect 3743 35581 3755 35584
rect 3697 35575 3755 35581
rect 4154 35572 4160 35584
rect 4212 35572 4218 35624
rect 2501 35547 2559 35553
rect 2501 35513 2513 35547
rect 2547 35544 2559 35547
rect 8846 35544 8852 35556
rect 2547 35516 8852 35544
rect 2547 35513 2559 35516
rect 2501 35507 2559 35513
rect 8846 35504 8852 35516
rect 8904 35504 8910 35556
rect 4982 35436 4988 35488
rect 5040 35476 5046 35488
rect 5350 35476 5356 35488
rect 5040 35448 5356 35476
rect 5040 35436 5046 35448
rect 5350 35436 5356 35448
rect 5408 35436 5414 35488
rect 10042 35476 10048 35488
rect 10003 35448 10048 35476
rect 10042 35436 10048 35448
rect 10100 35436 10106 35488
rect 1104 35386 10856 35408
rect 1104 35334 2582 35386
rect 2634 35334 2646 35386
rect 2698 35334 2710 35386
rect 2762 35334 2774 35386
rect 2826 35334 2838 35386
rect 2890 35334 5845 35386
rect 5897 35334 5909 35386
rect 5961 35334 5973 35386
rect 6025 35334 6037 35386
rect 6089 35334 6101 35386
rect 6153 35334 9109 35386
rect 9161 35334 9173 35386
rect 9225 35334 9237 35386
rect 9289 35334 9301 35386
rect 9353 35334 9365 35386
rect 9417 35334 10856 35386
rect 1104 35312 10856 35334
rect 3237 35275 3295 35281
rect 3237 35241 3249 35275
rect 3283 35272 3295 35275
rect 9766 35272 9772 35284
rect 3283 35244 9772 35272
rect 3283 35241 3295 35244
rect 3237 35235 3295 35241
rect 9766 35232 9772 35244
rect 9824 35232 9830 35284
rect 2501 35207 2559 35213
rect 2501 35173 2513 35207
rect 2547 35204 2559 35207
rect 8386 35204 8392 35216
rect 2547 35176 8392 35204
rect 2547 35173 2559 35176
rect 2501 35167 2559 35173
rect 8386 35164 8392 35176
rect 8444 35164 8450 35216
rect 6270 35136 6276 35148
rect 1688 35108 6276 35136
rect 1688 35077 1716 35108
rect 6270 35096 6276 35108
rect 6328 35096 6334 35148
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35037 1731 35071
rect 1673 35031 1731 35037
rect 2225 35071 2283 35077
rect 2225 35037 2237 35071
rect 2271 35037 2283 35071
rect 2406 35068 2412 35080
rect 2367 35040 2412 35068
rect 2225 35031 2283 35037
rect 937 35003 995 35009
rect 937 34969 949 35003
rect 983 35000 995 35003
rect 2240 35000 2268 35031
rect 2406 35028 2412 35040
rect 2464 35028 2470 35080
rect 3053 35071 3111 35077
rect 3053 35068 3065 35071
rect 2746 35040 3065 35068
rect 2746 35000 2774 35040
rect 3053 35037 3065 35040
rect 3099 35037 3111 35071
rect 3053 35031 3111 35037
rect 3237 35071 3295 35077
rect 3237 35037 3249 35071
rect 3283 35068 3295 35071
rect 3418 35068 3424 35080
rect 3283 35040 3424 35068
rect 3283 35037 3295 35040
rect 3237 35031 3295 35037
rect 3418 35028 3424 35040
rect 3476 35068 3482 35080
rect 4154 35068 4160 35080
rect 3476 35040 4160 35068
rect 3476 35028 3482 35040
rect 4154 35028 4160 35040
rect 4212 35028 4218 35080
rect 9766 35028 9772 35080
rect 9824 35068 9830 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9824 35040 9873 35068
rect 9824 35028 9830 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 9861 35031 9919 35037
rect 983 34972 2774 35000
rect 983 34969 995 34972
rect 937 34963 995 34969
rect 1486 34932 1492 34944
rect 1447 34904 1492 34932
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 10042 34932 10048 34944
rect 10003 34904 10048 34932
rect 10042 34892 10048 34904
rect 10100 34892 10106 34944
rect 1104 34842 10856 34864
rect 1104 34790 4213 34842
rect 4265 34790 4277 34842
rect 4329 34790 4341 34842
rect 4393 34790 4405 34842
rect 4457 34790 4469 34842
rect 4521 34790 7477 34842
rect 7529 34790 7541 34842
rect 7593 34790 7605 34842
rect 7657 34790 7669 34842
rect 7721 34790 7733 34842
rect 7785 34790 10856 34842
rect 1104 34768 10856 34790
rect 1489 34731 1547 34737
rect 1489 34697 1501 34731
rect 1535 34728 1547 34731
rect 1578 34728 1584 34740
rect 1535 34700 1584 34728
rect 1535 34697 1547 34700
rect 1489 34691 1547 34697
rect 1578 34688 1584 34700
rect 1636 34688 1642 34740
rect 2593 34663 2651 34669
rect 2593 34629 2605 34663
rect 2639 34660 2651 34663
rect 8662 34660 8668 34672
rect 2639 34632 8668 34660
rect 2639 34629 2651 34632
rect 2593 34623 2651 34629
rect 8662 34620 8668 34632
rect 8720 34620 8726 34672
rect 1578 34592 1584 34604
rect 1539 34564 1584 34592
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 2222 34592 2228 34604
rect 2183 34564 2228 34592
rect 2222 34552 2228 34564
rect 2280 34552 2286 34604
rect 2406 34592 2412 34604
rect 2367 34564 2412 34592
rect 2406 34552 2412 34564
rect 2464 34552 2470 34604
rect 3053 34595 3111 34601
rect 3053 34561 3065 34595
rect 3099 34592 3111 34595
rect 3234 34592 3240 34604
rect 3099 34564 3240 34592
rect 3099 34561 3111 34564
rect 3053 34555 3111 34561
rect 3234 34552 3240 34564
rect 3292 34552 3298 34604
rect 3234 34388 3240 34400
rect 3195 34360 3240 34388
rect 3234 34348 3240 34360
rect 3292 34348 3298 34400
rect 1104 34298 10856 34320
rect 1104 34246 2582 34298
rect 2634 34246 2646 34298
rect 2698 34246 2710 34298
rect 2762 34246 2774 34298
rect 2826 34246 2838 34298
rect 2890 34246 5845 34298
rect 5897 34246 5909 34298
rect 5961 34246 5973 34298
rect 6025 34246 6037 34298
rect 6089 34246 6101 34298
rect 6153 34246 9109 34298
rect 9161 34246 9173 34298
rect 9225 34246 9237 34298
rect 9289 34246 9301 34298
rect 9353 34246 9365 34298
rect 9417 34246 10856 34298
rect 1104 34224 10856 34246
rect 1762 34144 1768 34196
rect 1820 34184 1826 34196
rect 2222 34184 2228 34196
rect 1820 34156 2228 34184
rect 1820 34144 1826 34156
rect 2222 34144 2228 34156
rect 2280 34184 2286 34196
rect 3605 34187 3663 34193
rect 3605 34184 3617 34187
rect 2280 34156 3617 34184
rect 2280 34144 2286 34156
rect 3605 34153 3617 34156
rect 3651 34153 3663 34187
rect 3605 34147 3663 34153
rect 3973 34187 4031 34193
rect 3973 34153 3985 34187
rect 4019 34184 4031 34187
rect 9858 34184 9864 34196
rect 4019 34156 9864 34184
rect 4019 34153 4031 34156
rect 3973 34147 4031 34153
rect 9858 34144 9864 34156
rect 9916 34144 9922 34196
rect 3050 34116 3056 34128
rect 3011 34088 3056 34116
rect 3050 34076 3056 34088
rect 3108 34076 3114 34128
rect 11425 34051 11483 34057
rect 11425 34048 11437 34051
rect 1688 34020 11437 34048
rect 1688 33989 1716 34020
rect 11425 34017 11437 34020
rect 11471 34017 11483 34051
rect 11425 34011 11483 34017
rect 1673 33983 1731 33989
rect 1673 33949 1685 33983
rect 1719 33949 1731 33983
rect 1673 33943 1731 33949
rect 1946 33940 1952 33992
rect 2004 33980 2010 33992
rect 2133 33983 2191 33989
rect 2133 33980 2145 33983
rect 2004 33952 2145 33980
rect 2004 33940 2010 33952
rect 2133 33949 2145 33952
rect 2179 33949 2191 33983
rect 2133 33943 2191 33949
rect 2869 33983 2927 33989
rect 2869 33949 2881 33983
rect 2915 33980 2927 33983
rect 3326 33980 3332 33992
rect 2915 33952 3332 33980
rect 2915 33949 2927 33952
rect 2869 33943 2927 33949
rect 3326 33940 3332 33952
rect 3384 33940 3390 33992
rect 3605 33983 3663 33989
rect 3605 33949 3617 33983
rect 3651 33980 3663 33983
rect 3789 33983 3847 33989
rect 3789 33980 3801 33983
rect 3651 33952 3801 33980
rect 3651 33949 3663 33952
rect 3605 33943 3663 33949
rect 3789 33949 3801 33952
rect 3835 33949 3847 33983
rect 3789 33943 3847 33949
rect 3973 33983 4031 33989
rect 3973 33949 3985 33983
rect 4019 33949 4031 33983
rect 3973 33943 4031 33949
rect 3418 33872 3424 33924
rect 3476 33912 3482 33924
rect 3988 33912 4016 33943
rect 9674 33940 9680 33992
rect 9732 33980 9738 33992
rect 9861 33983 9919 33989
rect 9861 33980 9873 33983
rect 9732 33952 9873 33980
rect 9732 33940 9738 33952
rect 9861 33949 9873 33952
rect 9907 33949 9919 33983
rect 9861 33943 9919 33949
rect 3476 33884 4016 33912
rect 3476 33872 3482 33884
rect 1486 33844 1492 33856
rect 1447 33816 1492 33844
rect 1486 33804 1492 33816
rect 1544 33804 1550 33856
rect 2314 33844 2320 33856
rect 2275 33816 2320 33844
rect 2314 33804 2320 33816
rect 2372 33804 2378 33856
rect 5350 33804 5356 33856
rect 5408 33844 5414 33856
rect 5534 33844 5540 33856
rect 5408 33816 5540 33844
rect 5408 33804 5414 33816
rect 5534 33804 5540 33816
rect 5592 33804 5598 33856
rect 10042 33844 10048 33856
rect 10003 33816 10048 33844
rect 10042 33804 10048 33816
rect 10100 33804 10106 33856
rect 1104 33754 10856 33776
rect 1104 33702 4213 33754
rect 4265 33702 4277 33754
rect 4329 33702 4341 33754
rect 4393 33702 4405 33754
rect 4457 33702 4469 33754
rect 4521 33702 7477 33754
rect 7529 33702 7541 33754
rect 7593 33702 7605 33754
rect 7657 33702 7669 33754
rect 7721 33702 7733 33754
rect 7785 33702 10856 33754
rect 1104 33680 10856 33702
rect 2501 33643 2559 33649
rect 2501 33609 2513 33643
rect 2547 33640 2559 33643
rect 3145 33643 3203 33649
rect 2547 33612 2774 33640
rect 2547 33609 2559 33612
rect 2501 33603 2559 33609
rect 2746 33572 2774 33612
rect 3145 33609 3157 33643
rect 3191 33640 3203 33643
rect 9766 33640 9772 33652
rect 3191 33612 9772 33640
rect 3191 33609 3203 33612
rect 3145 33603 3203 33609
rect 9766 33600 9772 33612
rect 9824 33600 9830 33652
rect 1688 33544 2544 33572
rect 2746 33544 3556 33572
rect 1688 33513 1716 33544
rect 2516 33516 2544 33544
rect 1673 33507 1731 33513
rect 1673 33473 1685 33507
rect 1719 33473 1731 33507
rect 1673 33467 1731 33473
rect 1946 33464 1952 33516
rect 2004 33504 2010 33516
rect 2317 33507 2375 33513
rect 2317 33504 2329 33507
rect 2004 33476 2329 33504
rect 2004 33464 2010 33476
rect 2317 33473 2329 33476
rect 2363 33504 2375 33507
rect 2406 33504 2412 33516
rect 2363 33476 2412 33504
rect 2363 33473 2375 33476
rect 2317 33467 2375 33473
rect 2406 33464 2412 33476
rect 2464 33464 2470 33516
rect 2498 33464 2504 33516
rect 2556 33464 2562 33516
rect 2593 33507 2651 33513
rect 2593 33473 2605 33507
rect 2639 33504 2651 33507
rect 3053 33507 3111 33513
rect 3053 33504 3065 33507
rect 2639 33476 3065 33504
rect 2639 33473 2651 33476
rect 2593 33467 2651 33473
rect 2222 33396 2228 33448
rect 2280 33436 2286 33448
rect 2746 33436 2774 33476
rect 3053 33473 3065 33476
rect 3099 33473 3111 33507
rect 3053 33467 3111 33473
rect 3237 33507 3295 33513
rect 3237 33473 3249 33507
rect 3283 33504 3295 33507
rect 3418 33504 3424 33516
rect 3283 33476 3424 33504
rect 3283 33473 3295 33476
rect 3237 33467 3295 33473
rect 3418 33464 3424 33476
rect 3476 33464 3482 33516
rect 3528 33504 3556 33544
rect 7098 33504 7104 33516
rect 3528 33476 7104 33504
rect 7098 33464 7104 33476
rect 7156 33464 7162 33516
rect 9858 33504 9864 33516
rect 9819 33476 9864 33504
rect 9858 33464 9864 33476
rect 9916 33464 9922 33516
rect 2280 33408 2774 33436
rect 2280 33396 2286 33408
rect 1394 33260 1400 33312
rect 1452 33300 1458 33312
rect 1489 33303 1547 33309
rect 1489 33300 1501 33303
rect 1452 33272 1501 33300
rect 1452 33260 1458 33272
rect 1489 33269 1501 33272
rect 1535 33269 1547 33303
rect 10042 33300 10048 33312
rect 10003 33272 10048 33300
rect 1489 33263 1547 33269
rect 10042 33260 10048 33272
rect 10100 33260 10106 33312
rect 1104 33210 10856 33232
rect 1104 33158 2582 33210
rect 2634 33158 2646 33210
rect 2698 33158 2710 33210
rect 2762 33158 2774 33210
rect 2826 33158 2838 33210
rect 2890 33158 5845 33210
rect 5897 33158 5909 33210
rect 5961 33158 5973 33210
rect 6025 33158 6037 33210
rect 6089 33158 6101 33210
rect 6153 33158 9109 33210
rect 9161 33158 9173 33210
rect 9225 33158 9237 33210
rect 9289 33158 9301 33210
rect 9353 33158 9365 33210
rect 9417 33158 10856 33210
rect 1104 33136 10856 33158
rect 2869 33099 2927 33105
rect 2869 33065 2881 33099
rect 2915 33096 2927 33099
rect 2958 33096 2964 33108
rect 2915 33068 2964 33096
rect 2915 33065 2927 33068
rect 2869 33059 2927 33065
rect 2958 33056 2964 33068
rect 3016 33056 3022 33108
rect 3789 33099 3847 33105
rect 3789 33065 3801 33099
rect 3835 33096 3847 33099
rect 4798 33096 4804 33108
rect 3835 33068 4804 33096
rect 3835 33065 3847 33068
rect 3789 33059 3847 33065
rect 4798 33056 4804 33068
rect 4856 33056 4862 33108
rect 2314 32920 2320 32972
rect 2372 32960 2378 32972
rect 2498 32960 2504 32972
rect 2372 32932 2504 32960
rect 2372 32920 2378 32932
rect 2498 32920 2504 32932
rect 2556 32960 2562 32972
rect 4798 32960 4804 32972
rect 2556 32932 2774 32960
rect 2556 32920 2562 32932
rect 1210 32852 1216 32904
rect 1268 32892 1274 32904
rect 1673 32895 1731 32901
rect 1673 32892 1685 32895
rect 1268 32864 1685 32892
rect 1268 32852 1274 32864
rect 1673 32861 1685 32864
rect 1719 32861 1731 32895
rect 1673 32855 1731 32861
rect 2038 32852 2044 32904
rect 2096 32892 2102 32904
rect 2133 32895 2191 32901
rect 2133 32892 2145 32895
rect 2096 32864 2145 32892
rect 2096 32852 2102 32864
rect 2133 32861 2145 32864
rect 2179 32861 2191 32895
rect 2746 32892 2774 32932
rect 3068 32932 4804 32960
rect 3068 32901 3096 32932
rect 4798 32920 4804 32932
rect 4856 32920 4862 32972
rect 2869 32895 2927 32901
rect 2869 32892 2881 32895
rect 2746 32864 2881 32892
rect 2133 32855 2191 32861
rect 2869 32861 2881 32864
rect 2915 32861 2927 32895
rect 2869 32855 2927 32861
rect 3053 32895 3111 32901
rect 3053 32861 3065 32895
rect 3099 32861 3111 32895
rect 3053 32855 3111 32861
rect 3789 32895 3847 32901
rect 3789 32861 3801 32895
rect 3835 32861 3847 32895
rect 3789 32855 3847 32861
rect 3973 32895 4031 32901
rect 3973 32861 3985 32895
rect 4019 32892 4031 32895
rect 5534 32892 5540 32904
rect 4019 32864 5540 32892
rect 4019 32861 4031 32864
rect 3973 32855 4031 32861
rect 2884 32824 2912 32855
rect 3804 32824 3832 32855
rect 5534 32852 5540 32864
rect 5592 32852 5598 32904
rect 2884 32796 3832 32824
rect 1210 32716 1216 32768
rect 1268 32756 1274 32768
rect 1489 32759 1547 32765
rect 1489 32756 1501 32759
rect 1268 32728 1501 32756
rect 1268 32716 1274 32728
rect 1489 32725 1501 32728
rect 1535 32725 1547 32759
rect 2314 32756 2320 32768
rect 2275 32728 2320 32756
rect 1489 32719 1547 32725
rect 2314 32716 2320 32728
rect 2372 32716 2378 32768
rect 1104 32666 10856 32688
rect 1104 32614 4213 32666
rect 4265 32614 4277 32666
rect 4329 32614 4341 32666
rect 4393 32614 4405 32666
rect 4457 32614 4469 32666
rect 4521 32614 7477 32666
rect 7529 32614 7541 32666
rect 7593 32614 7605 32666
rect 7657 32614 7669 32666
rect 7721 32614 7733 32666
rect 7785 32614 10856 32666
rect 1104 32592 10856 32614
rect 1302 32512 1308 32564
rect 1360 32552 1366 32564
rect 1489 32555 1547 32561
rect 1489 32552 1501 32555
rect 1360 32524 1501 32552
rect 1360 32512 1366 32524
rect 1489 32521 1501 32524
rect 1535 32521 1547 32555
rect 2498 32552 2504 32564
rect 1489 32515 1547 32521
rect 1596 32524 2504 32552
rect 1302 32376 1308 32428
rect 1360 32416 1366 32428
rect 1596 32425 1624 32524
rect 2498 32512 2504 32524
rect 2556 32512 2562 32564
rect 3329 32555 3387 32561
rect 3329 32521 3341 32555
rect 3375 32552 3387 32555
rect 9674 32552 9680 32564
rect 3375 32524 9680 32552
rect 3375 32521 3387 32524
rect 3329 32515 3387 32521
rect 9674 32512 9680 32524
rect 9732 32512 9738 32564
rect 1946 32444 1952 32496
rect 2004 32484 2010 32496
rect 2409 32487 2467 32493
rect 2004 32456 2268 32484
rect 2004 32444 2010 32456
rect 1397 32419 1455 32425
rect 1397 32416 1409 32419
rect 1360 32388 1409 32416
rect 1360 32376 1366 32388
rect 1397 32385 1409 32388
rect 1443 32385 1455 32419
rect 1397 32379 1455 32385
rect 1581 32419 1639 32425
rect 1581 32385 1593 32419
rect 1627 32385 1639 32419
rect 2130 32416 2136 32428
rect 2091 32388 2136 32416
rect 1581 32379 1639 32385
rect 2130 32376 2136 32388
rect 2188 32376 2194 32428
rect 2240 32425 2268 32456
rect 2409 32453 2421 32487
rect 2455 32484 2467 32487
rect 6546 32484 6552 32496
rect 2455 32456 6552 32484
rect 2455 32453 2467 32456
rect 2409 32447 2467 32453
rect 6546 32444 6552 32456
rect 6604 32444 6610 32496
rect 2225 32419 2283 32425
rect 2225 32385 2237 32419
rect 2271 32385 2283 32419
rect 3237 32419 3295 32425
rect 3237 32416 3249 32419
rect 2225 32379 2283 32385
rect 2746 32388 3249 32416
rect 2148 32348 2176 32376
rect 2746 32348 2774 32388
rect 3237 32385 3249 32388
rect 3283 32385 3295 32419
rect 3237 32379 3295 32385
rect 3418 32376 3424 32428
rect 3476 32416 3482 32428
rect 3970 32416 3976 32428
rect 3476 32388 3976 32416
rect 3476 32376 3482 32388
rect 3970 32376 3976 32388
rect 4028 32376 4034 32428
rect 9861 32419 9919 32425
rect 9861 32385 9873 32419
rect 9907 32416 9919 32419
rect 11241 32419 11299 32425
rect 11241 32416 11253 32419
rect 9907 32388 11253 32416
rect 9907 32385 9919 32388
rect 9861 32379 9919 32385
rect 11241 32385 11253 32388
rect 11287 32385 11299 32419
rect 11241 32379 11299 32385
rect 2148 32320 2774 32348
rect 10042 32280 10048 32292
rect 10003 32252 10048 32280
rect 10042 32240 10048 32252
rect 10100 32240 10106 32292
rect 1486 32172 1492 32224
rect 1544 32212 1550 32224
rect 2314 32212 2320 32224
rect 1544 32184 2320 32212
rect 1544 32172 1550 32184
rect 2314 32172 2320 32184
rect 2372 32172 2378 32224
rect 1104 32122 10856 32144
rect 1104 32070 2582 32122
rect 2634 32070 2646 32122
rect 2698 32070 2710 32122
rect 2762 32070 2774 32122
rect 2826 32070 2838 32122
rect 2890 32070 5845 32122
rect 5897 32070 5909 32122
rect 5961 32070 5973 32122
rect 6025 32070 6037 32122
rect 6089 32070 6101 32122
rect 6153 32070 9109 32122
rect 9161 32070 9173 32122
rect 9225 32070 9237 32122
rect 9289 32070 9301 32122
rect 9353 32070 9365 32122
rect 9417 32070 10856 32122
rect 1104 32048 10856 32070
rect 1486 31968 1492 32020
rect 1544 32008 1550 32020
rect 1581 32011 1639 32017
rect 1581 32008 1593 32011
rect 1544 31980 1593 32008
rect 1544 31968 1550 31980
rect 1581 31977 1593 31980
rect 1627 31977 1639 32011
rect 3973 32011 4031 32017
rect 1581 31971 1639 31977
rect 2240 31980 2774 32008
rect 2240 31813 2268 31980
rect 2746 31940 2774 31980
rect 3973 31977 3985 32011
rect 4019 32008 4031 32011
rect 9858 32008 9864 32020
rect 4019 31980 9864 32008
rect 4019 31977 4031 31980
rect 3973 31971 4031 31977
rect 9858 31968 9864 31980
rect 9916 31968 9922 32020
rect 11517 31943 11575 31949
rect 11517 31940 11529 31943
rect 2746 31912 11529 31940
rect 11517 31909 11529 31912
rect 11563 31909 11575 31943
rect 11517 31903 11575 31909
rect 2314 31832 2320 31884
rect 2372 31872 2378 31884
rect 2372 31844 3832 31872
rect 2372 31832 2378 31844
rect 1765 31807 1823 31813
rect 1765 31773 1777 31807
rect 1811 31804 1823 31807
rect 2225 31807 2283 31813
rect 1811 31776 2176 31804
rect 1811 31773 1823 31776
rect 1765 31767 1823 31773
rect 2148 31736 2176 31776
rect 2225 31773 2237 31807
rect 2271 31773 2283 31807
rect 3418 31804 3424 31816
rect 2225 31767 2283 31773
rect 2332 31776 3424 31804
rect 2332 31736 2360 31776
rect 3418 31764 3424 31776
rect 3476 31764 3482 31816
rect 3804 31813 3832 31844
rect 3789 31807 3847 31813
rect 3789 31773 3801 31807
rect 3835 31773 3847 31807
rect 3970 31804 3976 31816
rect 3931 31776 3976 31804
rect 3789 31767 3847 31773
rect 3970 31764 3976 31776
rect 4028 31764 4034 31816
rect 4062 31764 4068 31816
rect 4120 31804 4126 31816
rect 7190 31804 7196 31816
rect 4120 31776 7196 31804
rect 4120 31764 4126 31776
rect 7190 31764 7196 31776
rect 7248 31764 7254 31816
rect 9861 31807 9919 31813
rect 9861 31773 9873 31807
rect 9907 31804 9919 31807
rect 11149 31807 11207 31813
rect 11149 31804 11161 31807
rect 9907 31776 11161 31804
rect 9907 31773 9919 31776
rect 9861 31767 9919 31773
rect 11149 31773 11161 31776
rect 11195 31773 11207 31807
rect 11149 31767 11207 31773
rect 2148 31708 2360 31736
rect 3602 31696 3608 31748
rect 3660 31696 3666 31748
rect 2406 31668 2412 31680
rect 2367 31640 2412 31668
rect 2406 31628 2412 31640
rect 2464 31628 2470 31680
rect 3620 31668 3648 31696
rect 3970 31668 3976 31680
rect 3620 31640 3976 31668
rect 3970 31628 3976 31640
rect 4028 31628 4034 31680
rect 10042 31668 10048 31680
rect 10003 31640 10048 31668
rect 10042 31628 10048 31640
rect 10100 31628 10106 31680
rect 1104 31578 10856 31600
rect 1104 31526 4213 31578
rect 4265 31526 4277 31578
rect 4329 31526 4341 31578
rect 4393 31526 4405 31578
rect 4457 31526 4469 31578
rect 4521 31526 7477 31578
rect 7529 31526 7541 31578
rect 7593 31526 7605 31578
rect 7657 31526 7669 31578
rect 7721 31526 7733 31578
rect 7785 31526 10856 31578
rect 1104 31504 10856 31526
rect 934 31356 940 31408
rect 992 31396 998 31408
rect 1489 31399 1547 31405
rect 1489 31396 1501 31399
rect 992 31368 1501 31396
rect 992 31356 998 31368
rect 1489 31365 1501 31368
rect 1535 31365 1547 31399
rect 10965 31399 11023 31405
rect 10965 31396 10977 31399
rect 1489 31359 1547 31365
rect 2746 31368 10977 31396
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31297 1823 31331
rect 1765 31291 1823 31297
rect 2225 31331 2283 31337
rect 2225 31297 2237 31331
rect 2271 31328 2283 31331
rect 2746 31328 2774 31368
rect 10965 31365 10977 31368
rect 11011 31365 11023 31399
rect 10965 31359 11023 31365
rect 2271 31300 2774 31328
rect 9861 31331 9919 31337
rect 2271 31297 2283 31300
rect 2225 31291 2283 31297
rect 9861 31297 9873 31331
rect 9907 31328 9919 31331
rect 11057 31331 11115 31337
rect 11057 31328 11069 31331
rect 9907 31300 11069 31328
rect 9907 31297 9919 31300
rect 9861 31291 9919 31297
rect 11057 31297 11069 31300
rect 11103 31297 11115 31331
rect 11057 31291 11115 31297
rect 1780 31260 1808 31291
rect 3050 31260 3056 31272
rect 1780 31232 3056 31260
rect 3050 31220 3056 31232
rect 3108 31220 3114 31272
rect 2406 31124 2412 31136
rect 2367 31096 2412 31124
rect 2406 31084 2412 31096
rect 2464 31084 2470 31136
rect 10042 31124 10048 31136
rect 10003 31096 10048 31124
rect 10042 31084 10048 31096
rect 10100 31084 10106 31136
rect 1104 31034 10856 31056
rect 1104 30982 2582 31034
rect 2634 30982 2646 31034
rect 2698 30982 2710 31034
rect 2762 30982 2774 31034
rect 2826 30982 2838 31034
rect 2890 30982 5845 31034
rect 5897 30982 5909 31034
rect 5961 30982 5973 31034
rect 6025 30982 6037 31034
rect 6089 30982 6101 31034
rect 6153 30982 9109 31034
rect 9161 30982 9173 31034
rect 9225 30982 9237 31034
rect 9289 30982 9301 31034
rect 9353 30982 9365 31034
rect 9417 30982 10856 31034
rect 1104 30960 10856 30982
rect 290 30676 296 30728
rect 348 30716 354 30728
rect 1673 30719 1731 30725
rect 1673 30716 1685 30719
rect 348 30688 1685 30716
rect 348 30676 354 30688
rect 1673 30685 1685 30688
rect 1719 30685 1731 30719
rect 2314 30716 2320 30728
rect 2275 30688 2320 30716
rect 1673 30679 1731 30685
rect 2314 30676 2320 30688
rect 2372 30676 2378 30728
rect 10137 30719 10195 30725
rect 10137 30685 10149 30719
rect 10183 30716 10195 30719
rect 10965 30719 11023 30725
rect 10965 30716 10977 30719
rect 10183 30688 10977 30716
rect 10183 30685 10195 30688
rect 10137 30679 10195 30685
rect 10965 30685 10977 30688
rect 11011 30685 11023 30719
rect 10965 30679 11023 30685
rect 1486 30580 1492 30592
rect 1447 30552 1492 30580
rect 1486 30540 1492 30552
rect 1544 30540 1550 30592
rect 1762 30540 1768 30592
rect 1820 30580 1826 30592
rect 2133 30583 2191 30589
rect 2133 30580 2145 30583
rect 1820 30552 2145 30580
rect 1820 30540 1826 30552
rect 2133 30549 2145 30552
rect 2179 30549 2191 30583
rect 2133 30543 2191 30549
rect 1104 30490 10856 30512
rect 1104 30438 4213 30490
rect 4265 30438 4277 30490
rect 4329 30438 4341 30490
rect 4393 30438 4405 30490
rect 4457 30438 4469 30490
rect 4521 30438 7477 30490
rect 7529 30438 7541 30490
rect 7593 30438 7605 30490
rect 7657 30438 7669 30490
rect 7721 30438 7733 30490
rect 7785 30438 10856 30490
rect 1104 30416 10856 30438
rect 1486 30336 1492 30388
rect 1544 30376 1550 30388
rect 1670 30376 1676 30388
rect 1544 30348 1676 30376
rect 1544 30336 1550 30348
rect 1670 30336 1676 30348
rect 1728 30336 1734 30388
rect 2130 30376 2136 30388
rect 1964 30348 2136 30376
rect 1581 30311 1639 30317
rect 1581 30277 1593 30311
rect 1627 30308 1639 30311
rect 1854 30308 1860 30320
rect 1627 30280 1860 30308
rect 1627 30277 1639 30280
rect 1581 30271 1639 30277
rect 1854 30268 1860 30280
rect 1912 30268 1918 30320
rect 1670 30240 1676 30252
rect 1631 30212 1676 30240
rect 1670 30200 1676 30212
rect 1728 30200 1734 30252
rect 1854 30132 1860 30184
rect 1912 30172 1918 30184
rect 1964 30172 1992 30348
rect 2130 30336 2136 30348
rect 2188 30336 2194 30388
rect 2130 30240 2136 30252
rect 2091 30212 2136 30240
rect 2130 30200 2136 30212
rect 2188 30200 2194 30252
rect 2958 30240 2964 30252
rect 2919 30212 2964 30240
rect 2958 30200 2964 30212
rect 3016 30200 3022 30252
rect 9858 30240 9864 30252
rect 9819 30212 9864 30240
rect 9858 30200 9864 30212
rect 9916 30200 9922 30252
rect 1912 30144 1992 30172
rect 1912 30132 1918 30144
rect 2038 30064 2044 30116
rect 2096 30104 2102 30116
rect 2317 30107 2375 30113
rect 2317 30104 2329 30107
rect 2096 30076 2329 30104
rect 2096 30064 2102 30076
rect 2317 30073 2329 30076
rect 2363 30073 2375 30107
rect 2317 30067 2375 30073
rect 1394 29996 1400 30048
rect 1452 30036 1458 30048
rect 2777 30039 2835 30045
rect 2777 30036 2789 30039
rect 1452 30008 2789 30036
rect 1452 29996 1458 30008
rect 2777 30005 2789 30008
rect 2823 30005 2835 30039
rect 10042 30036 10048 30048
rect 10003 30008 10048 30036
rect 2777 29999 2835 30005
rect 10042 29996 10048 30008
rect 10100 29996 10106 30048
rect 1104 29946 10856 29968
rect 1104 29894 2582 29946
rect 2634 29894 2646 29946
rect 2698 29894 2710 29946
rect 2762 29894 2774 29946
rect 2826 29894 2838 29946
rect 2890 29894 5845 29946
rect 5897 29894 5909 29946
rect 5961 29894 5973 29946
rect 6025 29894 6037 29946
rect 6089 29894 6101 29946
rect 6153 29894 9109 29946
rect 9161 29894 9173 29946
rect 9225 29894 9237 29946
rect 9289 29894 9301 29946
rect 9353 29894 9365 29946
rect 9417 29894 10856 29946
rect 1104 29872 10856 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 1670 29792 1676 29844
rect 1728 29832 1734 29844
rect 2225 29835 2283 29841
rect 2225 29832 2237 29835
rect 1728 29804 2237 29832
rect 1728 29792 1734 29804
rect 2225 29801 2237 29804
rect 2271 29801 2283 29835
rect 2225 29795 2283 29801
rect 2869 29835 2927 29841
rect 2869 29801 2881 29835
rect 2915 29832 2927 29835
rect 3050 29832 3056 29844
rect 2915 29804 3056 29832
rect 2915 29801 2927 29804
rect 2869 29795 2927 29801
rect 3050 29792 3056 29804
rect 3108 29792 3114 29844
rect 937 29699 995 29705
rect 937 29665 949 29699
rect 983 29696 995 29699
rect 1578 29696 1584 29708
rect 983 29668 1584 29696
rect 983 29665 995 29668
rect 937 29659 995 29665
rect 1578 29656 1584 29668
rect 1636 29656 1642 29708
rect 1762 29628 1768 29640
rect 1723 29600 1768 29628
rect 1762 29588 1768 29600
rect 1820 29588 1826 29640
rect 2409 29631 2467 29637
rect 2409 29597 2421 29631
rect 2455 29628 2467 29631
rect 2958 29628 2964 29640
rect 2455 29600 2964 29628
rect 2455 29597 2467 29600
rect 2409 29591 2467 29597
rect 2958 29588 2964 29600
rect 3016 29588 3022 29640
rect 3050 29588 3056 29640
rect 3108 29628 3114 29640
rect 3108 29600 3153 29628
rect 3108 29588 3114 29600
rect 3234 29452 3240 29504
rect 3292 29492 3298 29504
rect 3694 29492 3700 29504
rect 3292 29464 3700 29492
rect 3292 29452 3298 29464
rect 3694 29452 3700 29464
rect 3752 29452 3758 29504
rect 1104 29402 10856 29424
rect 1104 29350 4213 29402
rect 4265 29350 4277 29402
rect 4329 29350 4341 29402
rect 4393 29350 4405 29402
rect 4457 29350 4469 29402
rect 4521 29350 7477 29402
rect 7529 29350 7541 29402
rect 7593 29350 7605 29402
rect 7657 29350 7669 29402
rect 7721 29350 7733 29402
rect 7785 29350 10856 29402
rect 1104 29328 10856 29350
rect 2038 29248 2044 29300
rect 2096 29288 2102 29300
rect 2406 29288 2412 29300
rect 2096 29260 2412 29288
rect 2096 29248 2102 29260
rect 2406 29248 2412 29260
rect 2464 29288 2470 29300
rect 2464 29260 3096 29288
rect 2464 29248 2470 29260
rect 2774 29220 2780 29232
rect 2056 29192 2780 29220
rect 2056 29161 2084 29192
rect 2774 29180 2780 29192
rect 2832 29180 2838 29232
rect 2041 29155 2099 29161
rect 2041 29121 2053 29155
rect 2087 29121 2099 29155
rect 2041 29115 2099 29121
rect 2225 29155 2283 29161
rect 2225 29121 2237 29155
rect 2271 29152 2283 29155
rect 2406 29152 2412 29164
rect 2271 29124 2412 29152
rect 2271 29121 2283 29124
rect 2225 29115 2283 29121
rect 2406 29112 2412 29124
rect 2464 29152 2470 29164
rect 3068 29161 3096 29260
rect 3418 29248 3424 29300
rect 3476 29288 3482 29300
rect 3605 29291 3663 29297
rect 3605 29288 3617 29291
rect 3476 29260 3617 29288
rect 3476 29248 3482 29260
rect 3605 29257 3617 29260
rect 3651 29257 3663 29291
rect 3605 29251 3663 29257
rect 10962 29220 10968 29232
rect 10923 29192 10968 29220
rect 10962 29180 10968 29192
rect 11020 29180 11026 29232
rect 2869 29155 2927 29161
rect 2869 29152 2881 29155
rect 2464 29124 2881 29152
rect 2464 29112 2470 29124
rect 2869 29121 2881 29124
rect 2915 29121 2927 29155
rect 2869 29115 2927 29121
rect 3053 29155 3111 29161
rect 3053 29121 3065 29155
rect 3099 29121 3111 29155
rect 3786 29152 3792 29164
rect 3747 29124 3792 29152
rect 3053 29115 3111 29121
rect 3786 29112 3792 29124
rect 3844 29112 3850 29164
rect 2317 29087 2375 29093
rect 2317 29053 2329 29087
rect 2363 29084 2375 29087
rect 8018 29084 8024 29096
rect 2363 29056 8024 29084
rect 2363 29053 2375 29056
rect 2317 29047 2375 29053
rect 8018 29044 8024 29056
rect 8076 29044 8082 29096
rect 2869 29019 2927 29025
rect 2869 28985 2881 29019
rect 2915 29016 2927 29019
rect 4062 29016 4068 29028
rect 2915 28988 4068 29016
rect 2915 28985 2927 28988
rect 2869 28979 2927 28985
rect 4062 28976 4068 28988
rect 4120 28976 4126 29028
rect 1394 28908 1400 28960
rect 1452 28948 1458 28960
rect 2958 28948 2964 28960
rect 1452 28920 2964 28948
rect 1452 28908 1458 28920
rect 2958 28908 2964 28920
rect 3016 28908 3022 28960
rect 3050 28908 3056 28960
rect 3108 28948 3114 28960
rect 3418 28948 3424 28960
rect 3108 28920 3424 28948
rect 3108 28908 3114 28920
rect 3418 28908 3424 28920
rect 3476 28908 3482 28960
rect 4890 28908 4896 28960
rect 4948 28948 4954 28960
rect 5074 28948 5080 28960
rect 4948 28920 5080 28948
rect 4948 28908 4954 28920
rect 5074 28908 5080 28920
rect 5132 28908 5138 28960
rect 10134 28948 10140 28960
rect 10095 28920 10140 28948
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 1104 28858 10856 28880
rect 1104 28806 2582 28858
rect 2634 28806 2646 28858
rect 2698 28806 2710 28858
rect 2762 28806 2774 28858
rect 2826 28806 2838 28858
rect 2890 28806 5845 28858
rect 5897 28806 5909 28858
rect 5961 28806 5973 28858
rect 6025 28806 6037 28858
rect 6089 28806 6101 28858
rect 6153 28806 9109 28858
rect 9161 28806 9173 28858
rect 9225 28806 9237 28858
rect 9289 28806 9301 28858
rect 9353 28806 9365 28858
rect 9417 28806 10856 28858
rect 1104 28784 10856 28806
rect 382 28704 388 28756
rect 440 28744 446 28756
rect 2593 28747 2651 28753
rect 2593 28744 2605 28747
rect 440 28716 2605 28744
rect 440 28704 446 28716
rect 2593 28713 2605 28716
rect 2639 28713 2651 28747
rect 2593 28707 2651 28713
rect 4614 28704 4620 28756
rect 4672 28744 4678 28756
rect 4890 28744 4896 28756
rect 4672 28716 4896 28744
rect 4672 28704 4678 28716
rect 4890 28704 4896 28716
rect 4948 28704 4954 28756
rect 2041 28679 2099 28685
rect 2041 28645 2053 28679
rect 2087 28676 2099 28679
rect 5442 28676 5448 28688
rect 2087 28648 5448 28676
rect 2087 28645 2099 28648
rect 2041 28639 2099 28645
rect 5442 28636 5448 28648
rect 5500 28636 5506 28688
rect 2041 28543 2099 28549
rect 2041 28509 2053 28543
rect 2087 28509 2099 28543
rect 2041 28503 2099 28509
rect 2056 28472 2084 28503
rect 2774 28500 2780 28552
rect 2832 28540 2838 28552
rect 3970 28540 3976 28552
rect 2832 28512 2877 28540
rect 3931 28512 3976 28540
rect 2832 28500 2838 28512
rect 3970 28500 3976 28512
rect 4028 28500 4034 28552
rect 4706 28472 4712 28484
rect 2056 28444 4712 28472
rect 4706 28432 4712 28444
rect 4764 28432 4770 28484
rect 2682 28364 2688 28416
rect 2740 28404 2746 28416
rect 3789 28407 3847 28413
rect 3789 28404 3801 28407
rect 2740 28376 3801 28404
rect 2740 28364 2746 28376
rect 3789 28373 3801 28376
rect 3835 28373 3847 28407
rect 3789 28367 3847 28373
rect 1104 28314 10856 28336
rect 1104 28262 4213 28314
rect 4265 28262 4277 28314
rect 4329 28262 4341 28314
rect 4393 28262 4405 28314
rect 4457 28262 4469 28314
rect 4521 28262 7477 28314
rect 7529 28262 7541 28314
rect 7593 28262 7605 28314
rect 7657 28262 7669 28314
rect 7721 28262 7733 28314
rect 7785 28262 10856 28314
rect 1104 28240 10856 28262
rect 2774 28160 2780 28212
rect 2832 28200 2838 28212
rect 3789 28203 3847 28209
rect 3789 28200 3801 28203
rect 2832 28172 3801 28200
rect 2832 28160 2838 28172
rect 3789 28169 3801 28172
rect 3835 28169 3847 28203
rect 3789 28163 3847 28169
rect 1486 28132 1492 28144
rect 1447 28104 1492 28132
rect 1486 28092 1492 28104
rect 1544 28092 1550 28144
rect 2682 28132 2688 28144
rect 1780 28104 2688 28132
rect 1780 28073 1808 28104
rect 2682 28092 2688 28104
rect 2740 28092 2746 28144
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28033 1823 28067
rect 2314 28064 2320 28076
rect 2275 28036 2320 28064
rect 1765 28027 1823 28033
rect 2314 28024 2320 28036
rect 2372 28024 2378 28076
rect 2406 28024 2412 28076
rect 2464 28064 2470 28076
rect 2501 28067 2559 28073
rect 2501 28064 2513 28067
rect 2464 28036 2513 28064
rect 2464 28024 2470 28036
rect 2501 28033 2513 28036
rect 2547 28033 2559 28067
rect 2501 28027 2559 28033
rect 3050 28024 3056 28076
rect 3108 28064 3114 28076
rect 3329 28067 3387 28073
rect 3329 28064 3341 28067
rect 3108 28036 3341 28064
rect 3108 28024 3114 28036
rect 3329 28033 3341 28036
rect 3375 28033 3387 28067
rect 3329 28027 3387 28033
rect 3418 28024 3424 28076
rect 3476 28064 3482 28076
rect 3973 28067 4031 28073
rect 3973 28064 3985 28067
rect 3476 28036 3985 28064
rect 3476 28024 3482 28036
rect 3973 28033 3985 28036
rect 4019 28033 4031 28067
rect 3973 28027 4031 28033
rect 2317 27931 2375 27937
rect 2317 27897 2329 27931
rect 2363 27928 2375 27931
rect 4614 27928 4620 27940
rect 2363 27900 4620 27928
rect 2363 27897 2375 27900
rect 2317 27891 2375 27897
rect 4614 27888 4620 27900
rect 4672 27888 4678 27940
rect 1946 27820 1952 27872
rect 2004 27860 2010 27872
rect 3145 27863 3203 27869
rect 3145 27860 3157 27863
rect 2004 27832 3157 27860
rect 2004 27820 2010 27832
rect 3145 27829 3157 27832
rect 3191 27829 3203 27863
rect 3145 27823 3203 27829
rect 1104 27770 10856 27792
rect 1104 27718 2582 27770
rect 2634 27718 2646 27770
rect 2698 27718 2710 27770
rect 2762 27718 2774 27770
rect 2826 27718 2838 27770
rect 2890 27718 5845 27770
rect 5897 27718 5909 27770
rect 5961 27718 5973 27770
rect 6025 27718 6037 27770
rect 6089 27718 6101 27770
rect 6153 27718 9109 27770
rect 9161 27718 9173 27770
rect 9225 27718 9237 27770
rect 9289 27718 9301 27770
rect 9353 27718 9365 27770
rect 9417 27718 10856 27770
rect 1104 27696 10856 27718
rect 2406 27616 2412 27668
rect 2464 27656 2470 27668
rect 3786 27656 3792 27668
rect 2464 27628 3792 27656
rect 2464 27616 2470 27628
rect 3786 27616 3792 27628
rect 3844 27616 3850 27668
rect 10134 27616 10140 27668
rect 10192 27616 10198 27668
rect 2317 27591 2375 27597
rect 2317 27557 2329 27591
rect 2363 27588 2375 27591
rect 3973 27591 4031 27597
rect 2363 27560 3924 27588
rect 2363 27557 2375 27560
rect 2317 27551 2375 27557
rect 2866 27480 2872 27532
rect 2924 27520 2930 27532
rect 3145 27523 3203 27529
rect 3145 27520 3157 27523
rect 2924 27492 3157 27520
rect 2924 27480 2930 27492
rect 3145 27489 3157 27492
rect 3191 27489 3203 27523
rect 3896 27520 3924 27560
rect 3973 27557 3985 27591
rect 4019 27588 4031 27591
rect 9858 27588 9864 27600
rect 4019 27560 9864 27588
rect 4019 27557 4031 27560
rect 3973 27551 4031 27557
rect 9858 27548 9864 27560
rect 9916 27548 9922 27600
rect 7374 27520 7380 27532
rect 3896 27492 7380 27520
rect 3145 27483 3203 27489
rect 7374 27480 7380 27492
rect 7432 27480 7438 27532
rect 10152 27529 10180 27616
rect 10137 27523 10195 27529
rect 10137 27489 10149 27523
rect 10183 27489 10195 27523
rect 10137 27483 10195 27489
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27412 1458 27464
rect 2130 27452 2136 27464
rect 2091 27424 2136 27452
rect 2130 27412 2136 27424
rect 2188 27412 2194 27464
rect 2314 27452 2320 27464
rect 2275 27424 2320 27452
rect 2314 27412 2320 27424
rect 2372 27412 2378 27464
rect 2590 27412 2596 27464
rect 2648 27452 2654 27464
rect 3053 27455 3111 27461
rect 3053 27452 3065 27455
rect 2648 27424 3065 27452
rect 2648 27412 2654 27424
rect 3053 27421 3065 27424
rect 3099 27421 3111 27455
rect 3053 27415 3111 27421
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 2774 27344 2780 27396
rect 2832 27384 2838 27396
rect 3252 27384 3280 27415
rect 3786 27412 3792 27464
rect 3844 27461 3850 27464
rect 3844 27452 3853 27461
rect 3844 27424 3889 27452
rect 3844 27415 3853 27424
rect 3844 27412 3850 27415
rect 3970 27412 3976 27464
rect 4028 27452 4034 27464
rect 4614 27452 4620 27464
rect 4028 27424 4620 27452
rect 4028 27412 4034 27424
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 2832 27356 3280 27384
rect 2832 27344 2838 27356
rect 6270 27344 6276 27396
rect 6328 27384 6334 27396
rect 11057 27387 11115 27393
rect 11057 27384 11069 27387
rect 6328 27356 11069 27384
rect 6328 27344 6334 27356
rect 11057 27353 11069 27356
rect 11103 27353 11115 27387
rect 11057 27347 11115 27353
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 1854 27316 1860 27328
rect 1627 27288 1860 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 1854 27276 1860 27288
rect 1912 27276 1918 27328
rect 2866 27276 2872 27328
rect 2924 27316 2930 27328
rect 5718 27316 5724 27328
rect 2924 27288 5724 27316
rect 2924 27276 2930 27288
rect 5718 27276 5724 27288
rect 5776 27276 5782 27328
rect 1104 27226 10856 27248
rect 1104 27174 4213 27226
rect 4265 27174 4277 27226
rect 4329 27174 4341 27226
rect 4393 27174 4405 27226
rect 4457 27174 4469 27226
rect 4521 27174 7477 27226
rect 7529 27174 7541 27226
rect 7593 27174 7605 27226
rect 7657 27174 7669 27226
rect 7721 27174 7733 27226
rect 7785 27174 10856 27226
rect 1104 27152 10856 27174
rect 2314 27072 2320 27124
rect 2372 27112 2378 27124
rect 2372 27084 2544 27112
rect 2372 27072 2378 27084
rect 658 27004 664 27056
rect 716 27044 722 27056
rect 1581 27047 1639 27053
rect 1581 27044 1593 27047
rect 716 27016 1593 27044
rect 716 27004 722 27016
rect 1581 27013 1593 27016
rect 1627 27013 1639 27047
rect 1581 27007 1639 27013
rect 2516 27044 2544 27084
rect 3510 27072 3516 27124
rect 3568 27112 3574 27124
rect 4062 27112 4068 27124
rect 3568 27084 4068 27112
rect 3568 27072 3574 27084
rect 4062 27072 4068 27084
rect 4120 27072 4126 27124
rect 4525 27115 4583 27121
rect 4525 27081 4537 27115
rect 4571 27112 4583 27115
rect 4706 27112 4712 27124
rect 4571 27084 4712 27112
rect 4571 27081 4583 27084
rect 4525 27075 4583 27081
rect 4706 27072 4712 27084
rect 4764 27072 4770 27124
rect 3145 27047 3203 27053
rect 3145 27044 3157 27047
rect 2516 27016 3157 27044
rect 1857 26979 1915 26985
rect 1857 26945 1869 26979
rect 1903 26976 1915 26979
rect 1946 26976 1952 26988
rect 1903 26948 1952 26976
rect 1903 26945 1915 26948
rect 1857 26939 1915 26945
rect 1946 26936 1952 26948
rect 2004 26936 2010 26988
rect 2516 26985 2544 27016
rect 3145 27013 3157 27016
rect 3191 27013 3203 27047
rect 3145 27007 3203 27013
rect 3973 27047 4031 27053
rect 3973 27013 3985 27047
rect 4019 27044 4031 27047
rect 11149 27047 11207 27053
rect 11149 27044 11161 27047
rect 4019 27016 11161 27044
rect 4019 27013 4031 27016
rect 3973 27007 4031 27013
rect 11149 27013 11161 27016
rect 11195 27013 11207 27047
rect 11149 27007 11207 27013
rect 2501 26979 2559 26985
rect 2501 26945 2513 26979
rect 2547 26945 2559 26979
rect 2501 26939 2559 26945
rect 2590 26936 2596 26988
rect 2648 26976 2654 26988
rect 2648 26948 2741 26976
rect 2648 26936 2654 26948
rect 3050 26936 3056 26988
rect 3108 26976 3114 26988
rect 3329 26979 3387 26985
rect 3329 26976 3341 26979
rect 3108 26948 3341 26976
rect 3108 26936 3114 26948
rect 3329 26945 3341 26948
rect 3375 26945 3387 26979
rect 3881 26979 3939 26985
rect 3881 26976 3893 26979
rect 3329 26939 3387 26945
rect 3620 26948 3893 26976
rect 2222 26868 2228 26920
rect 2280 26908 2286 26920
rect 2608 26908 2636 26936
rect 2280 26880 2636 26908
rect 2280 26868 2286 26880
rect 2409 26843 2467 26849
rect 2409 26809 2421 26843
rect 2455 26840 2467 26843
rect 2866 26840 2872 26852
rect 2455 26812 2872 26840
rect 2455 26809 2467 26812
rect 2409 26803 2467 26809
rect 2866 26800 2872 26812
rect 2924 26800 2930 26852
rect 3620 26784 3648 26948
rect 3881 26945 3893 26948
rect 3927 26945 3939 26979
rect 3881 26939 3939 26945
rect 4065 26979 4123 26985
rect 4065 26945 4077 26979
rect 4111 26976 4123 26979
rect 4614 26976 4620 26988
rect 4111 26948 4620 26976
rect 4111 26945 4123 26948
rect 4065 26939 4123 26945
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26945 4767 26979
rect 10134 26976 10140 26988
rect 10095 26948 10140 26976
rect 4709 26939 4767 26945
rect 3694 26868 3700 26920
rect 3752 26908 3758 26920
rect 4724 26908 4752 26939
rect 10134 26936 10140 26948
rect 10192 26936 10198 26988
rect 3752 26880 4752 26908
rect 3752 26868 3758 26880
rect 3602 26732 3608 26784
rect 3660 26732 3666 26784
rect 1104 26682 10856 26704
rect 1104 26630 2582 26682
rect 2634 26630 2646 26682
rect 2698 26630 2710 26682
rect 2762 26630 2774 26682
rect 2826 26630 2838 26682
rect 2890 26630 5845 26682
rect 5897 26630 5909 26682
rect 5961 26630 5973 26682
rect 6025 26630 6037 26682
rect 6089 26630 6101 26682
rect 6153 26630 9109 26682
rect 9161 26630 9173 26682
rect 9225 26630 9237 26682
rect 9289 26630 9301 26682
rect 9353 26630 9365 26682
rect 9417 26630 10856 26682
rect 1104 26608 10856 26630
rect 1946 26528 1952 26580
rect 2004 26568 2010 26580
rect 3789 26571 3847 26577
rect 3789 26568 3801 26571
rect 2004 26540 3801 26568
rect 2004 26528 2010 26540
rect 3789 26537 3801 26540
rect 3835 26537 3847 26571
rect 3789 26531 3847 26537
rect 2406 26460 2412 26512
rect 2464 26500 2470 26512
rect 2590 26500 2596 26512
rect 2464 26472 2596 26500
rect 2464 26460 2470 26472
rect 2590 26460 2596 26472
rect 2648 26460 2654 26512
rect 3145 26503 3203 26509
rect 3145 26469 3157 26503
rect 3191 26500 3203 26503
rect 11241 26503 11299 26509
rect 11241 26500 11253 26503
rect 3191 26472 11253 26500
rect 3191 26469 3203 26472
rect 3145 26463 3203 26469
rect 11241 26469 11253 26472
rect 11287 26469 11299 26503
rect 11241 26463 11299 26469
rect 1578 26392 1584 26444
rect 1636 26432 1642 26444
rect 1946 26432 1952 26444
rect 1636 26404 1952 26432
rect 1636 26392 1642 26404
rect 1946 26392 1952 26404
rect 2004 26392 2010 26444
rect 1210 26324 1216 26376
rect 1268 26364 1274 26376
rect 1397 26367 1455 26373
rect 1397 26364 1409 26367
rect 1268 26336 1409 26364
rect 1268 26324 1274 26336
rect 1397 26333 1409 26336
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 1486 26324 1492 26376
rect 1544 26364 1550 26376
rect 2041 26367 2099 26373
rect 2041 26364 2053 26367
rect 1544 26336 2053 26364
rect 1544 26324 1550 26336
rect 2041 26333 2053 26336
rect 2087 26333 2099 26367
rect 2041 26327 2099 26333
rect 2130 26324 2136 26376
rect 2188 26364 2194 26376
rect 2961 26367 3019 26373
rect 2961 26364 2973 26367
rect 2188 26336 2973 26364
rect 2188 26324 2194 26336
rect 2961 26333 2973 26336
rect 3007 26333 3019 26367
rect 2961 26327 3019 26333
rect 3145 26367 3203 26373
rect 3145 26333 3157 26367
rect 3191 26333 3203 26367
rect 3145 26327 3203 26333
rect 3160 26296 3188 26327
rect 3510 26324 3516 26376
rect 3568 26364 3574 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3568 26336 3985 26364
rect 3568 26324 3574 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4706 26296 4712 26308
rect 3160 26268 4712 26296
rect 4706 26256 4712 26268
rect 4764 26256 4770 26308
rect 1578 26228 1584 26240
rect 1539 26200 1584 26228
rect 1578 26188 1584 26200
rect 1636 26188 1642 26240
rect 2225 26231 2283 26237
rect 2225 26197 2237 26231
rect 2271 26228 2283 26231
rect 2314 26228 2320 26240
rect 2271 26200 2320 26228
rect 2271 26197 2283 26200
rect 2225 26191 2283 26197
rect 2314 26188 2320 26200
rect 2372 26188 2378 26240
rect 1104 26138 10856 26160
rect 1104 26086 4213 26138
rect 4265 26086 4277 26138
rect 4329 26086 4341 26138
rect 4393 26086 4405 26138
rect 4457 26086 4469 26138
rect 4521 26086 7477 26138
rect 7529 26086 7541 26138
rect 7593 26086 7605 26138
rect 7657 26086 7669 26138
rect 7721 26086 7733 26138
rect 7785 26086 10856 26138
rect 1104 26064 10856 26086
rect 2133 25959 2191 25965
rect 2133 25925 2145 25959
rect 2179 25956 2191 25959
rect 4890 25956 4896 25968
rect 2179 25928 4896 25956
rect 2179 25925 2191 25928
rect 2133 25919 2191 25925
rect 4890 25916 4896 25928
rect 4948 25916 4954 25968
rect 1854 25888 1860 25900
rect 1815 25860 1860 25888
rect 1854 25848 1860 25860
rect 1912 25848 1918 25900
rect 2777 25891 2835 25897
rect 2777 25857 2789 25891
rect 2823 25888 2835 25891
rect 2958 25888 2964 25900
rect 2823 25860 2964 25888
rect 2823 25857 2835 25860
rect 2777 25851 2835 25857
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 2590 25820 2596 25832
rect 1872 25792 2596 25820
rect 1872 25764 1900 25792
rect 2590 25780 2596 25792
rect 2648 25780 2654 25832
rect 1854 25712 1860 25764
rect 1912 25712 1918 25764
rect 2038 25644 2044 25696
rect 2096 25684 2102 25696
rect 2593 25687 2651 25693
rect 2593 25684 2605 25687
rect 2096 25656 2605 25684
rect 2096 25644 2102 25656
rect 2593 25653 2605 25656
rect 2639 25653 2651 25687
rect 2593 25647 2651 25653
rect 1104 25594 10856 25616
rect 1104 25542 2582 25594
rect 2634 25542 2646 25594
rect 2698 25542 2710 25594
rect 2762 25542 2774 25594
rect 2826 25542 2838 25594
rect 2890 25542 5845 25594
rect 5897 25542 5909 25594
rect 5961 25542 5973 25594
rect 6025 25542 6037 25594
rect 6089 25542 6101 25594
rect 6153 25542 9109 25594
rect 9161 25542 9173 25594
rect 9225 25542 9237 25594
rect 9289 25542 9301 25594
rect 9353 25542 9365 25594
rect 9417 25542 10856 25594
rect 1104 25520 10856 25542
rect 1118 25440 1124 25492
rect 1176 25480 1182 25492
rect 2317 25483 2375 25489
rect 2317 25480 2329 25483
rect 1176 25452 2329 25480
rect 1176 25440 1182 25452
rect 2317 25449 2329 25452
rect 2363 25449 2375 25483
rect 4982 25480 4988 25492
rect 2317 25443 2375 25449
rect 2746 25452 4988 25480
rect 1857 25415 1915 25421
rect 1857 25381 1869 25415
rect 1903 25412 1915 25415
rect 2746 25412 2774 25452
rect 4982 25440 4988 25452
rect 5040 25440 5046 25492
rect 10134 25480 10140 25492
rect 10095 25452 10140 25480
rect 10134 25440 10140 25452
rect 10192 25440 10198 25492
rect 1903 25384 2774 25412
rect 1903 25381 1915 25384
rect 1857 25375 1915 25381
rect 3234 25372 3240 25424
rect 3292 25412 3298 25424
rect 3510 25412 3516 25424
rect 3292 25384 3516 25412
rect 3292 25372 3298 25384
rect 3510 25372 3516 25384
rect 3568 25372 3574 25424
rect 1857 25279 1915 25285
rect 1857 25245 1869 25279
rect 1903 25276 1915 25279
rect 2038 25276 2044 25288
rect 1903 25248 2044 25276
rect 1903 25245 1915 25248
rect 1857 25239 1915 25245
rect 2038 25236 2044 25248
rect 2096 25236 2102 25288
rect 2314 25276 2320 25288
rect 2275 25248 2320 25276
rect 2314 25236 2320 25248
rect 2372 25236 2378 25288
rect 3234 25276 3240 25288
rect 3195 25248 3240 25276
rect 3234 25236 3240 25248
rect 3292 25236 3298 25288
rect 2866 25100 2872 25152
rect 2924 25140 2930 25152
rect 3053 25143 3111 25149
rect 3053 25140 3065 25143
rect 2924 25112 3065 25140
rect 2924 25100 2930 25112
rect 3053 25109 3065 25112
rect 3099 25109 3111 25143
rect 3053 25103 3111 25109
rect 1104 25050 10856 25072
rect 1104 24998 4213 25050
rect 4265 24998 4277 25050
rect 4329 24998 4341 25050
rect 4393 24998 4405 25050
rect 4457 24998 4469 25050
rect 4521 24998 7477 25050
rect 7529 24998 7541 25050
rect 7593 24998 7605 25050
rect 7657 24998 7669 25050
rect 7721 24998 7733 25050
rect 7785 24998 10856 25050
rect 1104 24976 10856 24998
rect 2314 24896 2320 24948
rect 2372 24936 2378 24948
rect 2590 24936 2596 24948
rect 2372 24908 2596 24936
rect 2372 24896 2378 24908
rect 2590 24896 2596 24908
rect 2648 24896 2654 24948
rect 3053 24871 3111 24877
rect 3053 24837 3065 24871
rect 3099 24868 3111 24871
rect 3326 24868 3332 24880
rect 3099 24840 3332 24868
rect 3099 24837 3111 24840
rect 3053 24831 3111 24837
rect 3326 24828 3332 24840
rect 3384 24828 3390 24880
rect 10226 24828 10232 24880
rect 10284 24828 10290 24880
rect 1397 24803 1455 24809
rect 1397 24769 1409 24803
rect 1443 24800 1455 24803
rect 1486 24800 1492 24812
rect 1443 24772 1492 24800
rect 1443 24769 1455 24772
rect 1397 24763 1455 24769
rect 1486 24760 1492 24772
rect 1544 24760 1550 24812
rect 2317 24803 2375 24809
rect 2317 24769 2329 24803
rect 2363 24800 2375 24803
rect 2866 24800 2872 24812
rect 2363 24772 2872 24800
rect 2363 24769 2375 24772
rect 2317 24763 2375 24769
rect 2866 24760 2872 24772
rect 2924 24760 2930 24812
rect 3421 24803 3479 24809
rect 3421 24769 3433 24803
rect 3467 24800 3479 24803
rect 4614 24800 4620 24812
rect 3467 24772 4620 24800
rect 3467 24769 3479 24772
rect 3421 24763 3479 24769
rect 566 24692 572 24744
rect 624 24732 630 24744
rect 3436 24732 3464 24763
rect 4614 24760 4620 24772
rect 4672 24760 4678 24812
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24800 10195 24803
rect 10244 24800 10272 24828
rect 10183 24772 10272 24800
rect 10183 24769 10195 24772
rect 10137 24763 10195 24769
rect 624 24704 3464 24732
rect 624 24692 630 24704
rect 1581 24667 1639 24673
rect 1581 24633 1593 24667
rect 1627 24664 1639 24667
rect 2958 24664 2964 24676
rect 1627 24636 2964 24664
rect 1627 24633 1639 24636
rect 1581 24627 1639 24633
rect 2958 24624 2964 24636
rect 3016 24624 3022 24676
rect 5166 24664 5172 24676
rect 3252 24636 5172 24664
rect 2317 24599 2375 24605
rect 2317 24565 2329 24599
rect 2363 24596 2375 24599
rect 3252 24596 3280 24636
rect 5166 24624 5172 24636
rect 5224 24624 5230 24676
rect 2363 24568 3280 24596
rect 2363 24565 2375 24568
rect 2317 24559 2375 24565
rect 1104 24506 10856 24528
rect 1104 24454 2582 24506
rect 2634 24454 2646 24506
rect 2698 24454 2710 24506
rect 2762 24454 2774 24506
rect 2826 24454 2838 24506
rect 2890 24454 5845 24506
rect 5897 24454 5909 24506
rect 5961 24454 5973 24506
rect 6025 24454 6037 24506
rect 6089 24454 6101 24506
rect 6153 24454 9109 24506
rect 9161 24454 9173 24506
rect 9225 24454 9237 24506
rect 9289 24454 9301 24506
rect 9353 24454 9365 24506
rect 9417 24454 10856 24506
rect 1104 24432 10856 24454
rect 2409 24395 2467 24401
rect 2409 24361 2421 24395
rect 2455 24392 2467 24395
rect 5074 24392 5080 24404
rect 2455 24364 5080 24392
rect 2455 24361 2467 24364
rect 2409 24355 2467 24361
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 10134 24392 10140 24404
rect 10095 24364 10140 24392
rect 10134 24352 10140 24364
rect 10192 24352 10198 24404
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 1578 24148 1584 24200
rect 1636 24188 1642 24200
rect 2225 24191 2283 24197
rect 2225 24188 2237 24191
rect 1636 24160 2237 24188
rect 1636 24148 1642 24160
rect 2225 24157 2237 24160
rect 2271 24157 2283 24191
rect 3142 24188 3148 24200
rect 3103 24160 3148 24188
rect 2225 24151 2283 24157
rect 3142 24148 3148 24160
rect 3200 24148 3206 24200
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 2130 24052 2136 24064
rect 1627 24024 2136 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 2130 24012 2136 24024
rect 2188 24012 2194 24064
rect 2498 24012 2504 24064
rect 2556 24052 2562 24064
rect 2961 24055 3019 24061
rect 2961 24052 2973 24055
rect 2556 24024 2973 24052
rect 2556 24012 2562 24024
rect 2961 24021 2973 24024
rect 3007 24021 3019 24055
rect 2961 24015 3019 24021
rect 1104 23962 10856 23984
rect 1104 23910 4213 23962
rect 4265 23910 4277 23962
rect 4329 23910 4341 23962
rect 4393 23910 4405 23962
rect 4457 23910 4469 23962
rect 4521 23910 7477 23962
rect 7529 23910 7541 23962
rect 7593 23910 7605 23962
rect 7657 23910 7669 23962
rect 7721 23910 7733 23962
rect 7785 23910 10856 23962
rect 1104 23888 10856 23910
rect 1026 23740 1032 23792
rect 1084 23780 1090 23792
rect 2225 23783 2283 23789
rect 2225 23780 2237 23783
rect 1084 23752 2237 23780
rect 1084 23740 1090 23752
rect 2225 23749 2237 23752
rect 2271 23749 2283 23783
rect 2225 23743 2283 23749
rect 1210 23672 1216 23724
rect 1268 23712 1274 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 1268 23684 1409 23712
rect 1268 23672 1274 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 2498 23712 2504 23724
rect 2459 23684 2504 23712
rect 1397 23675 1455 23681
rect 2498 23672 2504 23684
rect 2556 23672 2562 23724
rect 9858 23712 9864 23724
rect 9819 23684 9864 23712
rect 9858 23672 9864 23684
rect 9916 23672 9922 23724
rect 1578 23508 1584 23520
rect 1539 23480 1584 23508
rect 1578 23468 1584 23480
rect 1636 23468 1642 23520
rect 10042 23508 10048 23520
rect 10003 23480 10048 23508
rect 10042 23468 10048 23480
rect 10100 23468 10106 23520
rect 1104 23418 10856 23440
rect 1104 23366 2582 23418
rect 2634 23366 2646 23418
rect 2698 23366 2710 23418
rect 2762 23366 2774 23418
rect 2826 23366 2838 23418
rect 2890 23366 5845 23418
rect 5897 23366 5909 23418
rect 5961 23366 5973 23418
rect 6025 23366 6037 23418
rect 6089 23366 6101 23418
rect 6153 23366 9109 23418
rect 9161 23366 9173 23418
rect 9225 23366 9237 23418
rect 9289 23366 9301 23418
rect 9353 23366 9365 23418
rect 9417 23366 10856 23418
rect 1104 23344 10856 23366
rect 1581 23307 1639 23313
rect 1581 23273 1593 23307
rect 1627 23304 1639 23307
rect 2498 23304 2504 23316
rect 1627 23276 2504 23304
rect 1627 23273 1639 23276
rect 1581 23267 1639 23273
rect 2498 23264 2504 23276
rect 2556 23264 2562 23316
rect 3053 23307 3111 23313
rect 3053 23273 3065 23307
rect 3099 23304 3111 23307
rect 3786 23304 3792 23316
rect 3099 23276 3792 23304
rect 3099 23273 3111 23276
rect 3053 23267 3111 23273
rect 3786 23264 3792 23276
rect 3844 23264 3850 23316
rect 9493 23307 9551 23313
rect 9493 23273 9505 23307
rect 9539 23304 9551 23307
rect 9858 23304 9864 23316
rect 9539 23276 9864 23304
rect 9539 23273 9551 23276
rect 9493 23267 9551 23273
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 10134 23304 10140 23316
rect 10095 23276 10140 23304
rect 10134 23264 10140 23276
rect 10192 23264 10198 23316
rect 2317 23239 2375 23245
rect 2317 23205 2329 23239
rect 2363 23236 2375 23239
rect 3510 23236 3516 23248
rect 2363 23208 3516 23236
rect 2363 23205 2375 23208
rect 2317 23199 2375 23205
rect 3510 23196 3516 23208
rect 3568 23196 3574 23248
rect 1578 23100 1584 23112
rect 1539 23072 1584 23100
rect 1578 23060 1584 23072
rect 1636 23060 1642 23112
rect 2130 23100 2136 23112
rect 2091 23072 2136 23100
rect 2130 23060 2136 23072
rect 2188 23060 2194 23112
rect 2958 23100 2964 23112
rect 2919 23072 2964 23100
rect 2958 23060 2964 23072
rect 3016 23060 3022 23112
rect 3510 23060 3516 23112
rect 3568 23100 3574 23112
rect 9309 23103 9367 23109
rect 9309 23100 9321 23103
rect 3568 23072 9321 23100
rect 3568 23060 3574 23072
rect 9309 23069 9321 23072
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 1104 22874 10856 22896
rect 1104 22822 4213 22874
rect 4265 22822 4277 22874
rect 4329 22822 4341 22874
rect 4393 22822 4405 22874
rect 4457 22822 4469 22874
rect 4521 22822 7477 22874
rect 7529 22822 7541 22874
rect 7593 22822 7605 22874
rect 7657 22822 7669 22874
rect 7721 22822 7733 22874
rect 7785 22822 10856 22874
rect 1104 22800 10856 22822
rect 2409 22763 2467 22769
rect 2409 22729 2421 22763
rect 2455 22760 2467 22763
rect 5350 22760 5356 22772
rect 2455 22732 5356 22760
rect 2455 22729 2467 22732
rect 2409 22723 2467 22729
rect 5350 22720 5356 22732
rect 5408 22720 5414 22772
rect 3786 22692 3792 22704
rect 1872 22664 3792 22692
rect 1872 22633 1900 22664
rect 3786 22652 3792 22664
rect 3844 22652 3850 22704
rect 1857 22627 1915 22633
rect 1857 22593 1869 22627
rect 1903 22593 1915 22627
rect 1857 22587 1915 22593
rect 2501 22627 2559 22633
rect 2501 22593 2513 22627
rect 2547 22624 2559 22627
rect 3142 22624 3148 22636
rect 2547 22596 2774 22624
rect 3103 22596 3148 22624
rect 2547 22593 2559 22596
rect 2501 22587 2559 22593
rect 2746 22488 2774 22596
rect 3142 22584 3148 22596
rect 3200 22584 3206 22636
rect 9858 22624 9864 22636
rect 9819 22596 9864 22624
rect 9858 22584 9864 22596
rect 9916 22584 9922 22636
rect 2961 22491 3019 22497
rect 2961 22488 2973 22491
rect 2746 22460 2973 22488
rect 2961 22457 2973 22460
rect 3007 22457 3019 22491
rect 2961 22451 3019 22457
rect 1857 22423 1915 22429
rect 1857 22389 1869 22423
rect 1903 22420 1915 22423
rect 3970 22420 3976 22432
rect 1903 22392 3976 22420
rect 1903 22389 1915 22392
rect 1857 22383 1915 22389
rect 3970 22380 3976 22392
rect 4028 22380 4034 22432
rect 10042 22420 10048 22432
rect 10003 22392 10048 22420
rect 10042 22380 10048 22392
rect 10100 22380 10106 22432
rect 1104 22330 10856 22352
rect 1104 22278 2582 22330
rect 2634 22278 2646 22330
rect 2698 22278 2710 22330
rect 2762 22278 2774 22330
rect 2826 22278 2838 22330
rect 2890 22278 5845 22330
rect 5897 22278 5909 22330
rect 5961 22278 5973 22330
rect 6025 22278 6037 22330
rect 6089 22278 6101 22330
rect 6153 22278 9109 22330
rect 9161 22278 9173 22330
rect 9225 22278 9237 22330
rect 9289 22278 9301 22330
rect 9353 22278 9365 22330
rect 9417 22278 10856 22330
rect 1104 22256 10856 22278
rect 3786 22216 3792 22228
rect 3747 22188 3792 22216
rect 3786 22176 3792 22188
rect 3844 22176 3850 22228
rect 1949 22083 2007 22089
rect 1949 22049 1961 22083
rect 1995 22080 2007 22083
rect 3418 22080 3424 22092
rect 1995 22052 3424 22080
rect 1995 22049 2007 22052
rect 1949 22043 2007 22049
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 22012 2283 22015
rect 2866 22012 2872 22024
rect 2271 21984 2728 22012
rect 2827 21984 2872 22012
rect 2271 21981 2283 21984
rect 2225 21975 2283 21981
rect 2700 21885 2728 21984
rect 2866 21972 2872 21984
rect 2924 21972 2930 22024
rect 3970 22012 3976 22024
rect 3931 21984 3976 22012
rect 3970 21972 3976 21984
rect 4028 21972 4034 22024
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 22012 9919 22015
rect 9950 22012 9956 22024
rect 9907 21984 9956 22012
rect 9907 21981 9919 21984
rect 9861 21975 9919 21981
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 2685 21879 2743 21885
rect 2685 21845 2697 21879
rect 2731 21845 2743 21879
rect 10042 21876 10048 21888
rect 10003 21848 10048 21876
rect 2685 21839 2743 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 1104 21786 10856 21808
rect 1104 21734 4213 21786
rect 4265 21734 4277 21786
rect 4329 21734 4341 21786
rect 4393 21734 4405 21786
rect 4457 21734 4469 21786
rect 4521 21734 7477 21786
rect 7529 21734 7541 21786
rect 7593 21734 7605 21786
rect 7657 21734 7669 21786
rect 7721 21734 7733 21786
rect 7785 21734 10856 21786
rect 1104 21712 10856 21734
rect 1762 21632 1768 21684
rect 1820 21672 1826 21684
rect 1857 21675 1915 21681
rect 1857 21672 1869 21675
rect 1820 21644 1869 21672
rect 1820 21632 1826 21644
rect 1857 21641 1869 21644
rect 1903 21641 1915 21675
rect 1857 21635 1915 21641
rect 2130 21632 2136 21684
rect 2188 21672 2194 21684
rect 2314 21672 2320 21684
rect 2188 21644 2320 21672
rect 2188 21632 2194 21644
rect 2314 21632 2320 21644
rect 2372 21632 2378 21684
rect 3237 21607 3295 21613
rect 3237 21573 3249 21607
rect 3283 21604 3295 21607
rect 3326 21604 3332 21616
rect 3283 21576 3332 21604
rect 3283 21573 3295 21576
rect 3237 21567 3295 21573
rect 3326 21564 3332 21576
rect 3384 21564 3390 21616
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21536 2007 21539
rect 2314 21536 2320 21548
rect 1995 21508 2320 21536
rect 1995 21505 2007 21508
rect 1949 21499 2007 21505
rect 2314 21496 2320 21508
rect 2372 21496 2378 21548
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21505 2927 21539
rect 3878 21536 3884 21548
rect 3839 21508 3884 21536
rect 2869 21499 2927 21505
rect 1762 21428 1768 21480
rect 1820 21468 1826 21480
rect 2884 21468 2912 21499
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 1820 21440 2912 21468
rect 1820 21428 1826 21440
rect 2498 21400 2504 21412
rect 2459 21372 2504 21400
rect 2498 21360 2504 21372
rect 2556 21360 2562 21412
rect 3142 21292 3148 21344
rect 3200 21332 3206 21344
rect 3697 21335 3755 21341
rect 3697 21332 3709 21335
rect 3200 21304 3709 21332
rect 3200 21292 3206 21304
rect 3697 21301 3709 21304
rect 3743 21301 3755 21335
rect 3697 21295 3755 21301
rect 1104 21242 10856 21264
rect 1104 21190 2582 21242
rect 2634 21190 2646 21242
rect 2698 21190 2710 21242
rect 2762 21190 2774 21242
rect 2826 21190 2838 21242
rect 2890 21190 5845 21242
rect 5897 21190 5909 21242
rect 5961 21190 5973 21242
rect 6025 21190 6037 21242
rect 6089 21190 6101 21242
rect 6153 21190 9109 21242
rect 9161 21190 9173 21242
rect 9225 21190 9237 21242
rect 9289 21190 9301 21242
rect 9353 21190 9365 21242
rect 9417 21190 10856 21242
rect 1104 21168 10856 21190
rect 1946 21128 1952 21140
rect 1907 21100 1952 21128
rect 1946 21088 1952 21100
rect 2004 21088 2010 21140
rect 2314 21088 2320 21140
rect 2372 21128 2378 21140
rect 3789 21131 3847 21137
rect 3789 21128 3801 21131
rect 2372 21100 3801 21128
rect 2372 21088 2378 21100
rect 3789 21097 3801 21100
rect 3835 21097 3847 21131
rect 3789 21091 3847 21097
rect 2774 21020 2780 21072
rect 2832 21060 2838 21072
rect 2869 21063 2927 21069
rect 2869 21060 2881 21063
rect 2832 21032 2881 21060
rect 2832 21020 2838 21032
rect 2869 21029 2881 21032
rect 2915 21060 2927 21063
rect 5258 21060 5264 21072
rect 2915 21032 5264 21060
rect 2915 21029 2927 21032
rect 2869 21023 2927 21029
rect 5258 21020 5264 21032
rect 5316 21020 5322 21072
rect 2041 20927 2099 20933
rect 2041 20893 2053 20927
rect 2087 20924 2099 20927
rect 3694 20924 3700 20936
rect 2087 20896 3700 20924
rect 2087 20893 2099 20896
rect 2041 20887 2099 20893
rect 3694 20884 3700 20896
rect 3752 20884 3758 20936
rect 3970 20924 3976 20936
rect 3931 20896 3976 20924
rect 3970 20884 3976 20896
rect 4028 20884 4034 20936
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 9861 20927 9919 20933
rect 9861 20924 9873 20927
rect 9824 20896 9873 20924
rect 9824 20884 9830 20896
rect 9861 20893 9873 20896
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 2498 20856 2504 20868
rect 2459 20828 2504 20856
rect 2498 20816 2504 20828
rect 2556 20816 2562 20868
rect 2685 20859 2743 20865
rect 2685 20825 2697 20859
rect 2731 20825 2743 20859
rect 2685 20819 2743 20825
rect 1762 20748 1768 20800
rect 1820 20788 1826 20800
rect 1946 20788 1952 20800
rect 1820 20760 1952 20788
rect 1820 20748 1826 20760
rect 1946 20748 1952 20760
rect 2004 20788 2010 20800
rect 2700 20788 2728 20819
rect 2004 20760 2728 20788
rect 2004 20748 2010 20760
rect 2958 20748 2964 20800
rect 3016 20788 3022 20800
rect 3510 20788 3516 20800
rect 3016 20760 3516 20788
rect 3016 20748 3022 20760
rect 3510 20748 3516 20760
rect 3568 20748 3574 20800
rect 10042 20788 10048 20800
rect 10003 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 1104 20698 10856 20720
rect 1104 20646 4213 20698
rect 4265 20646 4277 20698
rect 4329 20646 4341 20698
rect 4393 20646 4405 20698
rect 4457 20646 4469 20698
rect 4521 20646 7477 20698
rect 7529 20646 7541 20698
rect 7593 20646 7605 20698
rect 7657 20646 7669 20698
rect 7721 20646 7733 20698
rect 7785 20646 10856 20698
rect 1104 20624 10856 20646
rect 1581 20587 1639 20593
rect 1581 20553 1593 20587
rect 1627 20584 1639 20587
rect 1670 20584 1676 20596
rect 1627 20556 1676 20584
rect 1627 20553 1639 20556
rect 1581 20547 1639 20553
rect 1670 20544 1676 20556
rect 1728 20544 1734 20596
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 3050 20584 3056 20596
rect 2639 20556 3056 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 3050 20544 3056 20556
rect 3108 20544 3114 20596
rect 3694 20544 3700 20596
rect 3752 20584 3758 20596
rect 3881 20587 3939 20593
rect 3881 20584 3893 20587
rect 3752 20556 3893 20584
rect 3752 20544 3758 20556
rect 3881 20553 3893 20556
rect 3927 20553 3939 20587
rect 3881 20547 3939 20553
rect 4062 20544 4068 20596
rect 4120 20544 4126 20596
rect 9401 20587 9459 20593
rect 9401 20553 9413 20587
rect 9447 20584 9459 20587
rect 9858 20584 9864 20596
rect 9447 20556 9864 20584
rect 9447 20553 9459 20556
rect 9401 20547 9459 20553
rect 9858 20544 9864 20556
rect 9916 20544 9922 20596
rect 3510 20476 3516 20528
rect 3568 20516 3574 20528
rect 4080 20516 4108 20544
rect 3568 20488 4108 20516
rect 3568 20476 3574 20488
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 2314 20448 2320 20460
rect 1719 20420 2320 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 2314 20408 2320 20420
rect 2372 20408 2378 20460
rect 2774 20408 2780 20460
rect 2832 20448 2838 20460
rect 3418 20448 3424 20460
rect 2832 20420 2877 20448
rect 3379 20420 3424 20448
rect 2832 20408 2838 20420
rect 3418 20408 3424 20420
rect 3476 20408 3482 20460
rect 4062 20448 4068 20460
rect 4023 20420 4068 20448
rect 4062 20408 4068 20420
rect 4120 20408 4126 20460
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20417 9275 20451
rect 9858 20448 9864 20460
rect 9819 20420 9864 20448
rect 9217 20411 9275 20417
rect 3878 20340 3884 20392
rect 3936 20380 3942 20392
rect 9232 20380 9260 20411
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 3936 20352 9260 20380
rect 3936 20340 3942 20352
rect 3234 20244 3240 20256
rect 3195 20216 3240 20244
rect 3234 20204 3240 20216
rect 3292 20204 3298 20256
rect 10042 20244 10048 20256
rect 10003 20216 10048 20244
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 1104 20154 10856 20176
rect 1104 20102 2582 20154
rect 2634 20102 2646 20154
rect 2698 20102 2710 20154
rect 2762 20102 2774 20154
rect 2826 20102 2838 20154
rect 2890 20102 5845 20154
rect 5897 20102 5909 20154
rect 5961 20102 5973 20154
rect 6025 20102 6037 20154
rect 6089 20102 6101 20154
rect 6153 20102 9109 20154
rect 9161 20102 9173 20154
rect 9225 20102 9237 20154
rect 9289 20102 9301 20154
rect 9353 20102 9365 20154
rect 9417 20102 10856 20154
rect 1104 20080 10856 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2406 20040 2412 20052
rect 1995 20012 2412 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 3510 20040 3516 20052
rect 2639 20012 3516 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3234 19904 3240 19916
rect 2056 19876 3240 19904
rect 2056 19845 2084 19876
rect 3234 19864 3240 19876
rect 3292 19864 3298 19916
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19836 2743 19839
rect 3142 19836 3148 19848
rect 2731 19808 3148 19836
rect 2731 19805 2743 19808
rect 2685 19799 2743 19805
rect 3142 19796 3148 19808
rect 3200 19796 3206 19848
rect 9861 19839 9919 19845
rect 9861 19805 9873 19839
rect 9907 19836 9919 19839
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 9907 19808 10977 19836
rect 9907 19805 9919 19808
rect 9861 19799 9919 19805
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 4341 19771 4399 19777
rect 4341 19737 4353 19771
rect 4387 19768 4399 19771
rect 4614 19768 4620 19780
rect 4387 19740 4620 19768
rect 4387 19737 4399 19740
rect 4341 19731 4399 19737
rect 4614 19728 4620 19740
rect 4672 19728 4678 19780
rect 4249 19703 4307 19709
rect 4249 19669 4261 19703
rect 4295 19700 4307 19703
rect 4706 19700 4712 19712
rect 4295 19672 4712 19700
rect 4295 19669 4307 19672
rect 4249 19663 4307 19669
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 10042 19700 10048 19712
rect 10003 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 1104 19610 10856 19632
rect 1104 19558 4213 19610
rect 4265 19558 4277 19610
rect 4329 19558 4341 19610
rect 4393 19558 4405 19610
rect 4457 19558 4469 19610
rect 4521 19558 7477 19610
rect 7529 19558 7541 19610
rect 7593 19558 7605 19610
rect 7657 19558 7669 19610
rect 7721 19558 7733 19610
rect 7785 19558 10856 19610
rect 1104 19536 10856 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 2317 19499 2375 19505
rect 2317 19496 2329 19499
rect 2280 19468 2329 19496
rect 2280 19456 2286 19468
rect 2317 19465 2329 19468
rect 2363 19465 2375 19499
rect 2317 19459 2375 19465
rect 2406 19456 2412 19508
rect 2464 19496 2470 19508
rect 2869 19499 2927 19505
rect 2869 19496 2881 19499
rect 2464 19468 2881 19496
rect 2464 19456 2470 19468
rect 2869 19465 2881 19468
rect 2915 19465 2927 19499
rect 2869 19459 2927 19465
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 9950 19496 9956 19508
rect 3108 19468 3464 19496
rect 9911 19468 9956 19496
rect 3108 19456 3114 19468
rect 3436 19440 3464 19468
rect 9950 19456 9956 19468
rect 10008 19456 10014 19508
rect 3418 19388 3424 19440
rect 3476 19388 3482 19440
rect 1394 19360 1400 19372
rect 1355 19332 1400 19360
rect 1394 19320 1400 19332
rect 1452 19320 1458 19372
rect 2406 19360 2412 19372
rect 2367 19332 2412 19360
rect 2406 19320 2412 19332
rect 2464 19320 2470 19372
rect 3050 19360 3056 19372
rect 3011 19332 3056 19360
rect 3050 19320 3056 19332
rect 3108 19320 3114 19372
rect 10134 19360 10140 19372
rect 10095 19332 10140 19360
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 1104 19066 10856 19088
rect 1104 19014 2582 19066
rect 2634 19014 2646 19066
rect 2698 19014 2710 19066
rect 2762 19014 2774 19066
rect 2826 19014 2838 19066
rect 2890 19014 5845 19066
rect 5897 19014 5909 19066
rect 5961 19014 5973 19066
rect 6025 19014 6037 19066
rect 6089 19014 6101 19066
rect 6153 19014 9109 19066
rect 9161 19014 9173 19066
rect 9225 19014 9237 19066
rect 9289 19014 9301 19066
rect 9353 19014 9365 19066
rect 9417 19014 10856 19066
rect 1104 18992 10856 19014
rect 1857 18955 1915 18961
rect 1857 18921 1869 18955
rect 1903 18952 1915 18955
rect 2038 18952 2044 18964
rect 1903 18924 2044 18952
rect 1903 18921 1915 18924
rect 1857 18915 1915 18921
rect 2038 18912 2044 18924
rect 2096 18912 2102 18964
rect 9401 18955 9459 18961
rect 9401 18921 9413 18955
rect 9447 18952 9459 18955
rect 9766 18952 9772 18964
rect 9447 18924 9772 18952
rect 9447 18921 9459 18924
rect 9401 18915 9459 18921
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 3053 18887 3111 18893
rect 3053 18884 3065 18887
rect 2746 18856 3065 18884
rect 2746 18816 2774 18856
rect 3053 18853 3065 18856
rect 3099 18853 3111 18887
rect 3053 18847 3111 18853
rect 1964 18788 2774 18816
rect 1964 18757 1992 18788
rect 1949 18751 2007 18757
rect 1949 18717 1961 18751
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 2774 18748 2780 18760
rect 2639 18720 2780 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 2774 18708 2780 18720
rect 2832 18708 2838 18760
rect 3234 18748 3240 18760
rect 3195 18720 3240 18748
rect 3234 18708 3240 18720
rect 3292 18708 3298 18760
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9861 18751 9919 18757
rect 9861 18717 9873 18751
rect 9907 18748 9919 18751
rect 9950 18748 9956 18760
rect 9907 18720 9956 18748
rect 9907 18717 9919 18720
rect 9861 18711 9919 18717
rect 2314 18640 2320 18692
rect 2372 18680 2378 18692
rect 9232 18680 9260 18711
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 2372 18652 9260 18680
rect 2372 18640 2378 18652
rect 1946 18572 1952 18624
rect 2004 18612 2010 18624
rect 2409 18615 2467 18621
rect 2409 18612 2421 18615
rect 2004 18584 2421 18612
rect 2004 18572 2010 18584
rect 2409 18581 2421 18584
rect 2455 18581 2467 18615
rect 10042 18612 10048 18624
rect 10003 18584 10048 18612
rect 2409 18575 2467 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 1104 18522 10856 18544
rect 1104 18470 4213 18522
rect 4265 18470 4277 18522
rect 4329 18470 4341 18522
rect 4393 18470 4405 18522
rect 4457 18470 4469 18522
rect 4521 18470 7477 18522
rect 7529 18470 7541 18522
rect 7593 18470 7605 18522
rect 7657 18470 7669 18522
rect 7721 18470 7733 18522
rect 7785 18470 10856 18522
rect 1104 18448 10856 18470
rect 1854 18368 1860 18420
rect 1912 18408 1918 18420
rect 2133 18411 2191 18417
rect 2133 18408 2145 18411
rect 1912 18380 2145 18408
rect 1912 18368 1918 18380
rect 2133 18377 2145 18380
rect 2179 18377 2191 18411
rect 2133 18371 2191 18377
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 2685 18411 2743 18417
rect 2685 18408 2697 18411
rect 2464 18380 2697 18408
rect 2464 18368 2470 18380
rect 2685 18377 2697 18380
rect 2731 18377 2743 18411
rect 2685 18371 2743 18377
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 1946 18272 1952 18284
rect 1627 18244 1952 18272
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 3050 18272 3056 18284
rect 2915 18244 3056 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 9766 18232 9772 18284
rect 9824 18272 9830 18284
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9824 18244 9873 18272
rect 9824 18232 9830 18244
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 1489 18207 1547 18213
rect 1489 18173 1501 18207
rect 1535 18204 1547 18207
rect 2130 18204 2136 18216
rect 1535 18176 2136 18204
rect 1535 18173 1547 18176
rect 1489 18167 1547 18173
rect 2130 18164 2136 18176
rect 2188 18164 2194 18216
rect 10042 18068 10048 18080
rect 10003 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 1104 17978 10856 18000
rect 1104 17926 2582 17978
rect 2634 17926 2646 17978
rect 2698 17926 2710 17978
rect 2762 17926 2774 17978
rect 2826 17926 2838 17978
rect 2890 17926 5845 17978
rect 5897 17926 5909 17978
rect 5961 17926 5973 17978
rect 6025 17926 6037 17978
rect 6089 17926 6101 17978
rect 6153 17926 9109 17978
rect 9161 17926 9173 17978
rect 9225 17926 9237 17978
rect 9289 17926 9301 17978
rect 9353 17926 9365 17978
rect 9417 17926 10856 17978
rect 1104 17904 10856 17926
rect 1765 17867 1823 17873
rect 1765 17833 1777 17867
rect 1811 17864 1823 17867
rect 3602 17864 3608 17876
rect 1811 17836 3608 17864
rect 1811 17833 1823 17836
rect 1765 17827 1823 17833
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 9858 17864 9864 17876
rect 9819 17836 9864 17864
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17728 2927 17731
rect 2958 17728 2964 17740
rect 2915 17700 2964 17728
rect 2915 17697 2927 17700
rect 2869 17691 2927 17697
rect 2958 17688 2964 17700
rect 3016 17728 3022 17740
rect 3510 17728 3516 17740
rect 3016 17700 3516 17728
rect 3016 17688 3022 17700
rect 3510 17688 3516 17700
rect 3568 17688 3574 17740
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 1673 17663 1731 17669
rect 1673 17660 1685 17663
rect 1636 17632 1685 17660
rect 1636 17620 1642 17632
rect 1673 17629 1685 17632
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 2130 17620 2136 17672
rect 2188 17660 2194 17672
rect 2314 17660 2320 17672
rect 2188 17632 2320 17660
rect 2188 17620 2194 17632
rect 2314 17620 2320 17632
rect 2372 17660 2378 17672
rect 2501 17663 2559 17669
rect 2501 17660 2513 17663
rect 2372 17632 2513 17660
rect 2372 17620 2378 17632
rect 2501 17629 2513 17632
rect 2547 17629 2559 17663
rect 2501 17623 2559 17629
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 10045 17663 10103 17669
rect 10045 17660 10057 17663
rect 9732 17632 10057 17660
rect 9732 17620 9738 17632
rect 10045 17629 10057 17632
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 3878 17592 3884 17604
rect 2700 17564 3884 17592
rect 1946 17484 1952 17536
rect 2004 17524 2010 17536
rect 2590 17524 2596 17536
rect 2004 17496 2596 17524
rect 2004 17484 2010 17496
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 2700 17533 2728 17564
rect 3878 17552 3884 17564
rect 3936 17552 3942 17604
rect 2685 17527 2743 17533
rect 2685 17493 2697 17527
rect 2731 17493 2743 17527
rect 2685 17487 2743 17493
rect 2869 17527 2927 17533
rect 2869 17493 2881 17527
rect 2915 17524 2927 17527
rect 2958 17524 2964 17536
rect 2915 17496 2964 17524
rect 2915 17493 2927 17496
rect 2869 17487 2927 17493
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 1104 17434 10856 17456
rect 1104 17382 4213 17434
rect 4265 17382 4277 17434
rect 4329 17382 4341 17434
rect 4393 17382 4405 17434
rect 4457 17382 4469 17434
rect 4521 17382 7477 17434
rect 7529 17382 7541 17434
rect 7593 17382 7605 17434
rect 7657 17382 7669 17434
rect 7721 17382 7733 17434
rect 7785 17382 10856 17434
rect 1104 17360 10856 17382
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2685 17323 2743 17329
rect 2685 17320 2697 17323
rect 2280 17292 2697 17320
rect 2280 17280 2286 17292
rect 2685 17289 2697 17292
rect 2731 17289 2743 17323
rect 2685 17283 2743 17289
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 10134 17252 10140 17264
rect 2648 17224 10140 17252
rect 2648 17212 2654 17224
rect 10134 17212 10140 17224
rect 10192 17212 10198 17264
rect 1210 17144 1216 17196
rect 1268 17184 1274 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 1268 17156 1409 17184
rect 1268 17144 1274 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 2222 17184 2228 17196
rect 2183 17156 2228 17184
rect 1397 17147 1455 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 2866 17184 2872 17196
rect 2827 17156 2872 17184
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 9907 17156 11069 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 10042 17048 10048 17060
rect 10003 17020 10048 17048
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 1820 16952 2053 16980
rect 1820 16940 1826 16952
rect 2041 16949 2053 16952
rect 2087 16949 2099 16983
rect 2041 16943 2099 16949
rect 1104 16890 10856 16912
rect 1104 16838 2582 16890
rect 2634 16838 2646 16890
rect 2698 16838 2710 16890
rect 2762 16838 2774 16890
rect 2826 16838 2838 16890
rect 2890 16838 5845 16890
rect 5897 16838 5909 16890
rect 5961 16838 5973 16890
rect 6025 16838 6037 16890
rect 6089 16838 6101 16890
rect 6153 16838 9109 16890
rect 9161 16838 9173 16890
rect 9225 16838 9237 16890
rect 9289 16838 9301 16890
rect 9353 16838 9365 16890
rect 9417 16838 10856 16890
rect 1104 16816 10856 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 3142 16776 3148 16788
rect 3099 16748 3148 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 2958 16640 2964 16652
rect 2919 16612 2964 16640
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 1118 16532 1124 16584
rect 1176 16572 1182 16584
rect 1397 16575 1455 16581
rect 1397 16572 1409 16575
rect 1176 16544 1409 16572
rect 1176 16532 1182 16544
rect 1397 16541 1409 16544
rect 1443 16541 1455 16575
rect 1397 16535 1455 16541
rect 2777 16575 2835 16581
rect 2777 16541 2789 16575
rect 2823 16572 2835 16575
rect 9217 16575 9275 16581
rect 2823 16544 3004 16572
rect 2823 16541 2835 16544
rect 2777 16535 2835 16541
rect 2976 16516 3004 16544
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9858 16572 9864 16584
rect 9819 16544 9864 16572
rect 9217 16535 9275 16541
rect 2314 16464 2320 16516
rect 2372 16504 2378 16516
rect 2372 16476 2728 16504
rect 2372 16464 2378 16476
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 1581 16439 1639 16445
rect 1581 16436 1593 16439
rect 1452 16408 1593 16436
rect 1452 16396 1458 16408
rect 1581 16405 1593 16408
rect 1627 16405 1639 16439
rect 1581 16399 1639 16405
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 2593 16439 2651 16445
rect 2593 16436 2605 16439
rect 2556 16408 2605 16436
rect 2556 16396 2562 16408
rect 2593 16405 2605 16408
rect 2639 16405 2651 16439
rect 2700 16436 2728 16476
rect 2958 16464 2964 16516
rect 3016 16464 3022 16516
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 3108 16476 3153 16504
rect 3108 16464 3114 16476
rect 9232 16436 9260 16535
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 2700 16408 9260 16436
rect 9401 16439 9459 16445
rect 2593 16399 2651 16405
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9766 16436 9772 16448
rect 9447 16408 9772 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 1104 16346 10856 16368
rect 1104 16294 4213 16346
rect 4265 16294 4277 16346
rect 4329 16294 4341 16346
rect 4393 16294 4405 16346
rect 4457 16294 4469 16346
rect 4521 16294 7477 16346
rect 7529 16294 7541 16346
rect 7593 16294 7605 16346
rect 7657 16294 7669 16346
rect 7721 16294 7733 16346
rect 7785 16294 10856 16346
rect 1104 16272 10856 16294
rect 1949 16235 2007 16241
rect 1949 16201 1961 16235
rect 1995 16232 2007 16235
rect 2038 16232 2044 16244
rect 1995 16204 2044 16232
rect 1995 16201 2007 16204
rect 1949 16195 2007 16201
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 9401 16235 9459 16241
rect 9401 16201 9413 16235
rect 9447 16232 9459 16235
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 9447 16204 10977 16232
rect 9447 16201 9459 16204
rect 9401 16195 9459 16201
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 1486 16096 1492 16108
rect 1447 16068 1492 16096
rect 1486 16056 1492 16068
rect 1544 16056 1550 16108
rect 1762 16096 1768 16108
rect 1723 16068 1768 16096
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 2593 16099 2651 16105
rect 2593 16096 2605 16099
rect 1912 16068 2605 16096
rect 1912 16056 1918 16068
rect 2593 16065 2605 16068
rect 2639 16065 2651 16099
rect 3234 16096 3240 16108
rect 3195 16068 3240 16096
rect 2593 16059 2651 16065
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 4982 16056 4988 16108
rect 5040 16096 5046 16108
rect 9217 16099 9275 16105
rect 9217 16096 9229 16099
rect 5040 16068 9229 16096
rect 5040 16056 5046 16068
rect 9217 16065 9229 16068
rect 9263 16065 9275 16099
rect 9217 16059 9275 16065
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 11241 16099 11299 16105
rect 11241 16096 11253 16099
rect 9907 16068 11253 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 11241 16065 11253 16068
rect 11287 16065 11299 16099
rect 11241 16059 11299 16065
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 3053 15963 3111 15969
rect 3053 15960 3065 15963
rect 1780 15932 3065 15960
rect 1780 15901 1808 15932
rect 3053 15929 3065 15932
rect 3099 15929 3111 15963
rect 3053 15923 3111 15929
rect 1765 15895 1823 15901
rect 1765 15861 1777 15895
rect 1811 15861 1823 15895
rect 1765 15855 1823 15861
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 2096 15864 2421 15892
rect 2096 15852 2102 15864
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 10042 15892 10048 15904
rect 10003 15864 10048 15892
rect 2409 15855 2467 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 1104 15802 10856 15824
rect 1104 15750 2582 15802
rect 2634 15750 2646 15802
rect 2698 15750 2710 15802
rect 2762 15750 2774 15802
rect 2826 15750 2838 15802
rect 2890 15750 5845 15802
rect 5897 15750 5909 15802
rect 5961 15750 5973 15802
rect 6025 15750 6037 15802
rect 6089 15750 6101 15802
rect 6153 15750 9109 15802
rect 9161 15750 9173 15802
rect 9225 15750 9237 15802
rect 9289 15750 9301 15802
rect 9353 15750 9365 15802
rect 9417 15750 10856 15802
rect 1104 15728 10856 15750
rect 1489 15691 1547 15697
rect 1489 15657 1501 15691
rect 1535 15688 1547 15691
rect 1670 15688 1676 15700
rect 1535 15660 1676 15688
rect 1535 15657 1547 15660
rect 1489 15651 1547 15657
rect 1670 15648 1676 15660
rect 1728 15648 1734 15700
rect 2685 15691 2743 15697
rect 2685 15657 2697 15691
rect 2731 15688 2743 15691
rect 3050 15688 3056 15700
rect 2731 15660 3056 15688
rect 2731 15657 2743 15660
rect 2685 15651 2743 15657
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 2038 15552 2044 15564
rect 1412 15524 2044 15552
rect 1412 15493 1440 15524
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2314 15512 2320 15564
rect 2372 15512 2378 15564
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15552 2835 15555
rect 4062 15552 4068 15564
rect 2823 15524 4068 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 4062 15512 4068 15524
rect 4120 15552 4126 15564
rect 9674 15552 9680 15564
rect 4120 15524 9680 15552
rect 4120 15512 4126 15524
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15453 1455 15487
rect 1578 15484 1584 15496
rect 1539 15456 1584 15484
rect 1397 15447 1455 15453
rect 1578 15444 1584 15456
rect 1636 15444 1642 15496
rect 1762 15444 1768 15496
rect 1820 15484 1826 15496
rect 2332 15484 2360 15512
rect 2402 15487 2460 15493
rect 2402 15484 2414 15487
rect 1820 15456 2414 15484
rect 1820 15444 1826 15456
rect 2402 15453 2414 15456
rect 2448 15453 2460 15487
rect 2402 15447 2460 15453
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 10152 15416 10180 15447
rect 2516 15388 10180 15416
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 2516 15357 2544 15388
rect 2501 15351 2559 15357
rect 2501 15348 2513 15351
rect 2464 15320 2513 15348
rect 2464 15308 2470 15320
rect 2501 15317 2513 15320
rect 2547 15317 2559 15351
rect 2501 15311 2559 15317
rect 2590 15308 2596 15360
rect 2648 15348 2654 15360
rect 4982 15348 4988 15360
rect 2648 15320 4988 15348
rect 2648 15308 2654 15320
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 1104 15258 10856 15280
rect 1104 15206 4213 15258
rect 4265 15206 4277 15258
rect 4329 15206 4341 15258
rect 4393 15206 4405 15258
rect 4457 15206 4469 15258
rect 4521 15206 7477 15258
rect 7529 15206 7541 15258
rect 7593 15206 7605 15258
rect 7657 15206 7669 15258
rect 7721 15206 7733 15258
rect 7785 15206 10856 15258
rect 1104 15184 10856 15206
rect 1397 15147 1455 15153
rect 1397 15113 1409 15147
rect 1443 15144 1455 15147
rect 1486 15144 1492 15156
rect 1443 15116 1492 15144
rect 1443 15113 1455 15116
rect 1397 15107 1455 15113
rect 1486 15104 1492 15116
rect 1544 15104 1550 15156
rect 2593 15147 2651 15153
rect 2593 15113 2605 15147
rect 2639 15144 2651 15147
rect 2774 15144 2780 15156
rect 2639 15116 2780 15144
rect 2639 15113 2651 15116
rect 2593 15107 2651 15113
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 3234 15144 3240 15156
rect 2884 15116 3240 15144
rect 2884 15076 2912 15116
rect 3234 15104 3240 15116
rect 3292 15144 3298 15156
rect 3418 15144 3424 15156
rect 3292 15116 3424 15144
rect 3292 15104 3298 15116
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3602 15104 3608 15156
rect 3660 15144 3666 15156
rect 9030 15144 9036 15156
rect 3660 15116 9036 15144
rect 3660 15104 3666 15116
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9401 15147 9459 15153
rect 9401 15113 9413 15147
rect 9447 15144 9459 15147
rect 9858 15144 9864 15156
rect 9447 15116 9864 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 3513 15079 3571 15085
rect 2424 15048 2912 15076
rect 2976 15048 3464 15076
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 15008 1639 15011
rect 1627 14980 1808 15008
rect 1627 14977 1639 14980
rect 1581 14971 1639 14977
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 1673 14943 1731 14949
rect 1673 14940 1685 14943
rect 1452 14912 1685 14940
rect 1452 14900 1458 14912
rect 1673 14909 1685 14912
rect 1719 14909 1731 14943
rect 1780 14940 1808 14980
rect 1854 14968 1860 15020
rect 1912 15008 1918 15020
rect 1912 14980 1957 15008
rect 1912 14968 1918 14980
rect 2130 14968 2136 15020
rect 2188 15008 2194 15020
rect 2424 15017 2452 15048
rect 2409 15011 2467 15017
rect 2409 15008 2421 15011
rect 2188 14980 2421 15008
rect 2188 14968 2194 14980
rect 2409 14977 2421 14980
rect 2455 14977 2467 15011
rect 2409 14971 2467 14977
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 2976 15008 3004 15048
rect 2731 14980 3004 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 3050 14968 3056 15020
rect 3108 15008 3114 15020
rect 3145 15011 3203 15017
rect 3145 15008 3157 15011
rect 3108 14980 3157 15008
rect 3108 14968 3114 14980
rect 3145 14977 3157 14980
rect 3191 14977 3203 15011
rect 3145 14971 3203 14977
rect 3234 14968 3240 15020
rect 3292 15008 3298 15020
rect 3329 15011 3387 15017
rect 3329 15008 3341 15011
rect 3292 14980 3341 15008
rect 3292 14968 3298 14980
rect 3329 14977 3341 14980
rect 3375 14977 3387 15011
rect 3436 15008 3464 15048
rect 3513 15045 3525 15079
rect 3559 15076 3571 15079
rect 7926 15076 7932 15088
rect 3559 15048 7932 15076
rect 3559 15045 3571 15048
rect 3513 15039 3571 15045
rect 7926 15036 7932 15048
rect 7984 15036 7990 15088
rect 3602 15008 3608 15020
rect 3436 14980 3608 15008
rect 3329 14971 3387 14977
rect 3602 14968 3608 14980
rect 3660 14968 3666 15020
rect 9217 15011 9275 15017
rect 9217 14977 9229 15011
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 15008 9919 15011
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 9907 14980 11161 15008
rect 9907 14977 9919 14980
rect 9861 14971 9919 14977
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 3694 14940 3700 14952
rect 1780 14912 3700 14940
rect 1673 14903 1731 14909
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 3510 14832 3516 14884
rect 3568 14872 3574 14884
rect 9232 14872 9260 14971
rect 3568 14844 9260 14872
rect 3568 14832 3574 14844
rect 1857 14807 1915 14813
rect 1857 14773 1869 14807
rect 1903 14804 1915 14807
rect 3878 14804 3884 14816
rect 1903 14776 3884 14804
rect 1903 14773 1915 14776
rect 1857 14767 1915 14773
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 10042 14804 10048 14816
rect 10003 14776 10048 14804
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 1104 14714 10856 14736
rect 1104 14662 2582 14714
rect 2634 14662 2646 14714
rect 2698 14662 2710 14714
rect 2762 14662 2774 14714
rect 2826 14662 2838 14714
rect 2890 14662 5845 14714
rect 5897 14662 5909 14714
rect 5961 14662 5973 14714
rect 6025 14662 6037 14714
rect 6089 14662 6101 14714
rect 6153 14662 9109 14714
rect 9161 14662 9173 14714
rect 9225 14662 9237 14714
rect 9289 14662 9301 14714
rect 9353 14662 9365 14714
rect 9417 14662 10856 14714
rect 1104 14640 10856 14662
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 1912 14572 4445 14600
rect 1912 14560 1918 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 3752 14504 3801 14532
rect 3752 14492 3758 14504
rect 3789 14501 3801 14504
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 4706 14464 4712 14476
rect 3252 14436 4712 14464
rect 2130 14396 2136 14408
rect 2091 14368 2136 14396
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3252 14405 3280 14436
rect 4706 14424 4712 14436
rect 4764 14424 4770 14476
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3237 14359 3295 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4212 14368 4629 14396
rect 4212 14356 4218 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 9907 14368 10977 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 3145 14331 3203 14337
rect 2240 14300 2774 14328
rect 2240 14269 2268 14300
rect 2225 14263 2283 14269
rect 2225 14229 2237 14263
rect 2271 14229 2283 14263
rect 2746 14260 2774 14300
rect 3145 14297 3157 14331
rect 3191 14328 3203 14331
rect 11333 14331 11391 14337
rect 11333 14328 11345 14331
rect 3191 14300 11345 14328
rect 3191 14297 3203 14300
rect 3145 14291 3203 14297
rect 11333 14297 11345 14300
rect 11379 14297 11391 14331
rect 11333 14291 11391 14297
rect 8938 14260 8944 14272
rect 2746 14232 8944 14260
rect 2225 14223 2283 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 1104 14170 10856 14192
rect 1104 14118 4213 14170
rect 4265 14118 4277 14170
rect 4329 14118 4341 14170
rect 4393 14118 4405 14170
rect 4457 14118 4469 14170
rect 4521 14118 7477 14170
rect 7529 14118 7541 14170
rect 7593 14118 7605 14170
rect 7657 14118 7669 14170
rect 7721 14118 7733 14170
rect 7785 14118 10856 14170
rect 1104 14096 10856 14118
rect 2593 14059 2651 14065
rect 2593 14025 2605 14059
rect 2639 14056 2651 14059
rect 3050 14056 3056 14068
rect 2639 14028 3056 14056
rect 2639 14025 2651 14028
rect 2593 14019 2651 14025
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14025 3387 14059
rect 3329 14019 3387 14025
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 9858 14056 9864 14068
rect 4019 14028 9864 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 3344 13988 3372 14019
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 9766 13988 9772 14000
rect 2087 13960 2774 13988
rect 3344 13960 9772 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 1854 13920 1860 13932
rect 1815 13892 1860 13920
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2501 13923 2559 13929
rect 2501 13920 2513 13923
rect 2188 13892 2513 13920
rect 2188 13880 2194 13892
rect 2501 13889 2513 13892
rect 2547 13889 2559 13923
rect 2501 13883 2559 13889
rect 2746 13852 2774 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 3050 13880 3056 13932
rect 3108 13920 3114 13932
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 3108 13892 3157 13920
rect 3108 13880 3114 13892
rect 3145 13889 3157 13892
rect 3191 13920 3203 13923
rect 3326 13920 3332 13932
rect 3191 13892 3332 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3326 13880 3332 13892
rect 3384 13880 3390 13932
rect 3602 13880 3608 13932
rect 3660 13920 3666 13932
rect 3786 13920 3792 13932
rect 3660 13892 3792 13920
rect 3660 13880 3666 13892
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 4617 13923 4675 13929
rect 4617 13920 4629 13923
rect 4212 13892 4629 13920
rect 4212 13880 4218 13892
rect 4617 13889 4629 13892
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 3418 13852 3424 13864
rect 2746 13824 3424 13852
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 3936 13824 4476 13852
rect 3936 13812 3942 13824
rect 3142 13744 3148 13796
rect 3200 13784 3206 13796
rect 3326 13784 3332 13796
rect 3200 13756 3332 13784
rect 3200 13744 3206 13756
rect 3326 13744 3332 13756
rect 3384 13744 3390 13796
rect 4448 13793 4476 13824
rect 4433 13787 4491 13793
rect 4433 13753 4445 13787
rect 4479 13753 4491 13787
rect 4433 13747 4491 13753
rect 3418 13676 3424 13728
rect 3476 13716 3482 13728
rect 4062 13716 4068 13728
rect 3476 13688 4068 13716
rect 3476 13676 3482 13688
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 1104 13626 10856 13648
rect 1104 13574 2582 13626
rect 2634 13574 2646 13626
rect 2698 13574 2710 13626
rect 2762 13574 2774 13626
rect 2826 13574 2838 13626
rect 2890 13574 5845 13626
rect 5897 13574 5909 13626
rect 5961 13574 5973 13626
rect 6025 13574 6037 13626
rect 6089 13574 6101 13626
rect 6153 13574 9109 13626
rect 9161 13574 9173 13626
rect 9225 13574 9237 13626
rect 9289 13574 9301 13626
rect 9353 13574 9365 13626
rect 9417 13574 10856 13626
rect 1104 13552 10856 13574
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 2958 13512 2964 13524
rect 2915 13484 2964 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 2774 13404 2780 13456
rect 2832 13444 2838 13456
rect 3234 13444 3240 13456
rect 2832 13416 3240 13444
rect 2832 13404 2838 13416
rect 3234 13404 3240 13416
rect 3292 13404 3298 13456
rect 1673 13379 1731 13385
rect 1673 13345 1685 13379
rect 1719 13376 1731 13379
rect 1946 13376 1952 13388
rect 1719 13348 1952 13376
rect 1719 13345 1731 13348
rect 1673 13339 1731 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 3510 13376 3516 13388
rect 2792 13348 3516 13376
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 2792 13317 2820 13348
rect 3510 13336 3516 13348
rect 3568 13336 3574 13388
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13277 2835 13311
rect 2777 13271 2835 13277
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3142 13308 3148 13320
rect 3007 13280 3148 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 4341 13311 4399 13317
rect 4341 13277 4353 13311
rect 4387 13308 4399 13311
rect 4614 13308 4620 13320
rect 4387 13280 4620 13308
rect 4387 13277 4399 13280
rect 4341 13271 4399 13277
rect 4614 13268 4620 13280
rect 4672 13268 4678 13320
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 9950 13308 9956 13320
rect 9907 13280 9956 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 3234 13200 3240 13252
rect 3292 13240 3298 13252
rect 4157 13243 4215 13249
rect 4157 13240 4169 13243
rect 3292 13212 4169 13240
rect 3292 13200 3298 13212
rect 4157 13209 4169 13212
rect 4203 13209 4215 13243
rect 4157 13203 4215 13209
rect 10042 13172 10048 13184
rect 10003 13144 10048 13172
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 1104 13082 10856 13104
rect 1104 13030 4213 13082
rect 4265 13030 4277 13082
rect 4329 13030 4341 13082
rect 4393 13030 4405 13082
rect 4457 13030 4469 13082
rect 4521 13030 7477 13082
rect 7529 13030 7541 13082
rect 7593 13030 7605 13082
rect 7657 13030 7669 13082
rect 7721 13030 7733 13082
rect 7785 13030 10856 13082
rect 1104 13008 10856 13030
rect 9401 12971 9459 12977
rect 9401 12937 9413 12971
rect 9447 12968 9459 12971
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 9447 12940 11069 12968
rect 9447 12937 9459 12940
rect 9401 12931 9459 12937
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 11057 12931 11115 12937
rect 2958 12860 2964 12912
rect 3016 12860 3022 12912
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 2038 12832 2044 12844
rect 1719 12804 2044 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2976 12832 3004 12860
rect 3142 12832 3148 12844
rect 2976 12804 3148 12832
rect 3142 12792 3148 12804
rect 3200 12832 3206 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 3200 12804 9229 12832
rect 3200 12792 3206 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9858 12832 9864 12844
rect 9819 12804 9864 12832
rect 9217 12795 9275 12801
rect 9858 12792 9864 12804
rect 9916 12792 9922 12844
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1486 12764 1492 12776
rect 1443 12736 1492 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1486 12724 1492 12736
rect 1544 12724 1550 12776
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12764 2743 12767
rect 2774 12764 2780 12776
rect 2731 12736 2780 12764
rect 2731 12733 2743 12736
rect 2685 12727 2743 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 2924 12736 2973 12764
rect 2924 12724 2930 12736
rect 2961 12733 2973 12736
rect 3007 12733 3019 12767
rect 2961 12727 3019 12733
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 3510 12696 3516 12708
rect 3200 12668 3516 12696
rect 3200 12656 3206 12668
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 10042 12628 10048 12640
rect 10003 12600 10048 12628
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 1104 12538 10856 12560
rect 1104 12486 2582 12538
rect 2634 12486 2646 12538
rect 2698 12486 2710 12538
rect 2762 12486 2774 12538
rect 2826 12486 2838 12538
rect 2890 12486 5845 12538
rect 5897 12486 5909 12538
rect 5961 12486 5973 12538
rect 6025 12486 6037 12538
rect 6089 12486 6101 12538
rect 6153 12486 9109 12538
rect 9161 12486 9173 12538
rect 9225 12486 9237 12538
rect 9289 12486 9301 12538
rect 9353 12486 9365 12538
rect 9417 12486 10856 12538
rect 1104 12464 10856 12486
rect 2777 12427 2835 12433
rect 2777 12393 2789 12427
rect 2823 12424 2835 12427
rect 7834 12424 7840 12436
rect 2823 12396 7840 12424
rect 2823 12393 2835 12396
rect 2777 12387 2835 12393
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 1673 12291 1731 12297
rect 1673 12257 1685 12291
rect 1719 12288 1731 12291
rect 3418 12288 3424 12300
rect 1719 12260 3424 12288
rect 1719 12257 1731 12260
rect 1673 12251 1731 12257
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3878 12220 3884 12232
rect 3007 12192 3884 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9824 12192 9873 12220
rect 9824 12180 9830 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 1104 11994 10856 12016
rect 1104 11942 4213 11994
rect 4265 11942 4277 11994
rect 4329 11942 4341 11994
rect 4393 11942 4405 11994
rect 4457 11942 4469 11994
rect 4521 11942 7477 11994
rect 7529 11942 7541 11994
rect 7593 11942 7605 11994
rect 7657 11942 7669 11994
rect 7721 11942 7733 11994
rect 7785 11942 10856 11994
rect 1104 11920 10856 11942
rect 2777 11883 2835 11889
rect 2777 11849 2789 11883
rect 2823 11880 2835 11883
rect 6178 11880 6184 11892
rect 2823 11852 6184 11880
rect 2823 11849 2835 11852
rect 2777 11843 2835 11849
rect 6178 11840 6184 11852
rect 6236 11840 6242 11892
rect 9950 11880 9956 11892
rect 9911 11852 9956 11880
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 2222 11744 2228 11756
rect 1719 11716 2228 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3326 11744 3332 11756
rect 3007 11716 3332 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 10134 11744 10140 11756
rect 10095 11716 10140 11744
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 1397 11679 1455 11685
rect 1397 11676 1409 11679
rect 1360 11648 1409 11676
rect 1360 11636 1366 11648
rect 1397 11645 1409 11648
rect 1443 11645 1455 11679
rect 1397 11639 1455 11645
rect 1104 11450 10856 11472
rect 1104 11398 2582 11450
rect 2634 11398 2646 11450
rect 2698 11398 2710 11450
rect 2762 11398 2774 11450
rect 2826 11398 2838 11450
rect 2890 11398 5845 11450
rect 5897 11398 5909 11450
rect 5961 11398 5973 11450
rect 6025 11398 6037 11450
rect 6089 11398 6101 11450
rect 6153 11398 9109 11450
rect 9161 11398 9173 11450
rect 9225 11398 9237 11450
rect 9289 11398 9301 11450
rect 9353 11398 9365 11450
rect 9417 11398 10856 11450
rect 1104 11376 10856 11398
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 8202 11336 8208 11348
rect 2823 11308 8208 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 10965 11339 11023 11345
rect 10965 11336 10977 11339
rect 9447 11308 10977 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 10965 11305 10977 11308
rect 11011 11305 11023 11339
rect 10965 11299 11023 11305
rect 1578 11228 1584 11280
rect 1636 11268 1642 11280
rect 6730 11268 6736 11280
rect 1636 11240 6736 11268
rect 1636 11228 1642 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2406 11200 2412 11212
rect 1719 11172 2412 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 3510 11160 3516 11212
rect 3568 11200 3574 11212
rect 3568 11172 6914 11200
rect 3568 11160 3574 11172
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2924 11104 2973 11132
rect 2924 11092 2930 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11132 3847 11135
rect 3878 11132 3884 11144
rect 3835 11104 3884 11132
rect 3835 11101 3847 11104
rect 3789 11095 3847 11101
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 6886 11132 6914 11172
rect 9217 11135 9275 11141
rect 9217 11132 9229 11135
rect 6886 11104 9229 11132
rect 9217 11101 9229 11104
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11101 9919 11135
rect 9861 11095 9919 11101
rect 9876 11064 9904 11095
rect 3988 11036 9904 11064
rect 3988 11005 4016 11036
rect 3973 10999 4031 11005
rect 3973 10965 3985 10999
rect 4019 10965 4031 10999
rect 10042 10996 10048 11008
rect 10003 10968 10048 10996
rect 3973 10959 4031 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 1104 10906 10856 10928
rect 1104 10854 4213 10906
rect 4265 10854 4277 10906
rect 4329 10854 4341 10906
rect 4393 10854 4405 10906
rect 4457 10854 4469 10906
rect 4521 10854 7477 10906
rect 7529 10854 7541 10906
rect 7593 10854 7605 10906
rect 7657 10854 7669 10906
rect 7721 10854 7733 10906
rect 7785 10854 10856 10906
rect 1104 10832 10856 10854
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1762 10656 1768 10668
rect 1719 10628 1768 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1762 10616 1768 10628
rect 1820 10616 1826 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2866 10656 2872 10668
rect 2731 10628 2872 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2866 10616 2872 10628
rect 2924 10656 2930 10668
rect 3694 10656 3700 10668
rect 2924 10628 3700 10656
rect 2924 10616 2930 10628
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 9861 10659 9919 10665
rect 9861 10656 9873 10659
rect 6886 10628 9873 10656
rect 1302 10548 1308 10600
rect 1360 10588 1366 10600
rect 1397 10591 1455 10597
rect 1397 10588 1409 10591
rect 1360 10560 1409 10588
rect 1360 10548 1366 10560
rect 1397 10557 1409 10560
rect 1443 10557 1455 10591
rect 1397 10551 1455 10557
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 6886 10452 6914 10628
rect 9861 10625 9873 10628
rect 9907 10625 9919 10659
rect 9861 10619 9919 10625
rect 10042 10452 10048 10464
rect 2915 10424 6914 10452
rect 10003 10424 10048 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 1104 10362 10856 10384
rect 1104 10310 2582 10362
rect 2634 10310 2646 10362
rect 2698 10310 2710 10362
rect 2762 10310 2774 10362
rect 2826 10310 2838 10362
rect 2890 10310 5845 10362
rect 5897 10310 5909 10362
rect 5961 10310 5973 10362
rect 6025 10310 6037 10362
rect 6089 10310 6101 10362
rect 6153 10310 9109 10362
rect 9161 10310 9173 10362
rect 9225 10310 9237 10362
rect 9289 10310 9301 10362
rect 9353 10310 9365 10362
rect 9417 10310 10856 10362
rect 1104 10288 10856 10310
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 6638 10248 6644 10260
rect 2823 10220 6644 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 2958 10180 2964 10192
rect 1688 10152 2964 10180
rect 1688 10121 1716 10152
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 3142 10140 3148 10192
rect 3200 10140 3206 10192
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10081 1731 10115
rect 1673 10075 1731 10081
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 3160 10112 3188 10140
rect 2832 10084 3188 10112
rect 2832 10072 2838 10084
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3142 10044 3148 10056
rect 3007 10016 3148 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 1104 9818 10856 9840
rect 1104 9766 4213 9818
rect 4265 9766 4277 9818
rect 4329 9766 4341 9818
rect 4393 9766 4405 9818
rect 4457 9766 4469 9818
rect 4521 9766 7477 9818
rect 7529 9766 7541 9818
rect 7593 9766 7605 9818
rect 7657 9766 7669 9818
rect 7721 9766 7733 9818
rect 7785 9766 10856 9818
rect 1104 9744 10856 9766
rect 2777 9707 2835 9713
rect 2777 9673 2789 9707
rect 2823 9704 2835 9707
rect 3510 9704 3516 9716
rect 2823 9676 3516 9704
rect 2823 9673 2835 9676
rect 2777 9667 2835 9673
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 10134 9636 10140 9648
rect 2700 9608 10140 9636
rect 1762 9528 1768 9580
rect 1820 9568 1826 9580
rect 2700 9577 2728 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 1820 9540 2697 9568
rect 1820 9528 1826 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2899 9571 2957 9577
rect 2899 9537 2911 9571
rect 2945 9568 2957 9571
rect 4062 9568 4068 9580
rect 2945 9540 4068 9568
rect 2945 9537 2957 9540
rect 2899 9531 2957 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 8386 9528 8392 9580
rect 8444 9568 8450 9580
rect 9861 9571 9919 9577
rect 9861 9568 9873 9571
rect 8444 9540 9873 9568
rect 8444 9528 8450 9540
rect 9861 9537 9873 9540
rect 9907 9537 9919 9571
rect 9861 9531 9919 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2774 9500 2780 9512
rect 1719 9472 2780 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3970 9500 3976 9512
rect 3099 9472 3976 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 2961 9435 3019 9441
rect 2961 9401 2973 9435
rect 3007 9432 3019 9435
rect 3418 9432 3424 9444
rect 3007 9404 3424 9432
rect 3007 9401 3019 9404
rect 2961 9395 3019 9401
rect 3418 9392 3424 9404
rect 3476 9392 3482 9444
rect 10042 9432 10048 9444
rect 10003 9404 10048 9432
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 1104 9274 10856 9296
rect 1104 9222 2582 9274
rect 2634 9222 2646 9274
rect 2698 9222 2710 9274
rect 2762 9222 2774 9274
rect 2826 9222 2838 9274
rect 2890 9222 5845 9274
rect 5897 9222 5909 9274
rect 5961 9222 5973 9274
rect 6025 9222 6037 9274
rect 6089 9222 6101 9274
rect 6153 9222 9109 9274
rect 9161 9222 9173 9274
rect 9225 9222 9237 9274
rect 9289 9222 9301 9274
rect 9353 9222 9365 9274
rect 9417 9222 10856 9274
rect 1104 9200 10856 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3786 9160 3792 9172
rect 3476 9132 3792 9160
rect 3476 9120 3482 9132
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 9401 9163 9459 9169
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 11057 9163 11115 9169
rect 11057 9160 11069 9163
rect 9447 9132 11069 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 11057 9129 11069 9132
rect 11103 9129 11115 9163
rect 11057 9123 11115 9129
rect 2409 9095 2467 9101
rect 2409 9061 2421 9095
rect 2455 9092 2467 9095
rect 2455 9064 9904 9092
rect 2455 9061 2467 9064
rect 2409 9055 2467 9061
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 1811 8928 2237 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 3326 8956 3332 8968
rect 2915 8928 3332 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 2240 8888 2268 8919
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 3786 8956 3792 8968
rect 3747 8928 3792 8956
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 9876 8965 9904 9064
rect 9217 8959 9275 8965
rect 9217 8956 9229 8959
rect 4120 8928 9229 8956
rect 4120 8916 4126 8928
rect 9217 8925 9229 8928
rect 9263 8925 9275 8959
rect 9217 8919 9275 8925
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 2958 8888 2964 8900
rect 2240 8860 2964 8888
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 8386 8888 8392 8900
rect 3068 8860 8392 8888
rect 3068 8829 3096 8860
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 3053 8823 3111 8829
rect 3053 8789 3065 8823
rect 3099 8789 3111 8823
rect 3970 8820 3976 8832
rect 3883 8792 3976 8820
rect 3053 8783 3111 8789
rect 3970 8780 3976 8792
rect 4028 8820 4034 8832
rect 9214 8820 9220 8832
rect 4028 8792 9220 8820
rect 4028 8780 4034 8792
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 1104 8730 10856 8752
rect 1104 8678 4213 8730
rect 4265 8678 4277 8730
rect 4329 8678 4341 8730
rect 4393 8678 4405 8730
rect 4457 8678 4469 8730
rect 4521 8678 7477 8730
rect 7529 8678 7541 8730
rect 7593 8678 7605 8730
rect 7657 8678 7669 8730
rect 7721 8678 7733 8730
rect 7785 8678 10856 8730
rect 1104 8656 10856 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 4062 8616 4068 8628
rect 1627 8588 4068 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 9447 8588 11161 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8480 2559 8483
rect 3142 8480 3148 8492
rect 2547 8452 3148 8480
rect 2547 8449 2559 8452
rect 2501 8443 2559 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4062 8480 4068 8492
rect 3752 8452 4068 8480
rect 3752 8440 3758 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 9214 8480 9220 8492
rect 9175 8452 9220 8480
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 2685 8347 2743 8353
rect 2685 8313 2697 8347
rect 2731 8344 2743 8347
rect 9876 8344 9904 8443
rect 2731 8316 9904 8344
rect 2731 8313 2743 8316
rect 2685 8307 2743 8313
rect 10042 8276 10048 8288
rect 10003 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 1104 8186 10856 8208
rect 1104 8134 2582 8186
rect 2634 8134 2646 8186
rect 2698 8134 2710 8186
rect 2762 8134 2774 8186
rect 2826 8134 2838 8186
rect 2890 8134 5845 8186
rect 5897 8134 5909 8186
rect 5961 8134 5973 8186
rect 6025 8134 6037 8186
rect 6089 8134 6101 8186
rect 6153 8134 9109 8186
rect 9161 8134 9173 8186
rect 9225 8134 9237 8186
rect 9289 8134 9301 8186
rect 9353 8134 9365 8186
rect 9417 8134 10856 8186
rect 1104 8112 10856 8134
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1762 7936 1768 7948
rect 1719 7908 1768 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7837 3111 7871
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 3053 7831 3111 7837
rect 3068 7800 3096 7831
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 4798 7800 4804 7812
rect 3068 7772 4804 7800
rect 4798 7760 4804 7772
rect 4856 7760 4862 7812
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 9030 7732 9036 7744
rect 3191 7704 9036 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 1104 7642 10856 7664
rect 1104 7590 4213 7642
rect 4265 7590 4277 7642
rect 4329 7590 4341 7642
rect 4393 7590 4405 7642
rect 4457 7590 4469 7642
rect 4521 7590 7477 7642
rect 7529 7590 7541 7642
rect 7593 7590 7605 7642
rect 7657 7590 7669 7642
rect 7721 7590 7733 7642
rect 7785 7590 10856 7642
rect 1104 7568 10856 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3602 7528 3608 7540
rect 2915 7500 3608 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3602 7488 3608 7500
rect 3660 7488 3666 7540
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 3292 7432 3648 7460
rect 3292 7420 3298 7432
rect 1302 7352 1308 7404
rect 1360 7392 1366 7404
rect 1397 7395 1455 7401
rect 1397 7392 1409 7395
rect 1360 7364 1409 7392
rect 1360 7352 1366 7364
rect 1397 7361 1409 7364
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 2774 7392 2780 7404
rect 2731 7364 2780 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 3620 7401 3648 7432
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9732 7364 9873 7392
rect 9732 7352 9738 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 3510 7324 3516 7336
rect 1719 7296 3516 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 3602 7188 3608 7200
rect 3563 7160 3608 7188
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 10042 7188 10048 7200
rect 10003 7160 10048 7188
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 1104 7098 10856 7120
rect 1104 7046 2582 7098
rect 2634 7046 2646 7098
rect 2698 7046 2710 7098
rect 2762 7046 2774 7098
rect 2826 7046 2838 7098
rect 2890 7046 5845 7098
rect 5897 7046 5909 7098
rect 5961 7046 5973 7098
rect 6025 7046 6037 7098
rect 6089 7046 6101 7098
rect 6153 7046 9109 7098
rect 9161 7046 9173 7098
rect 9225 7046 9237 7098
rect 9289 7046 9301 7098
rect 9353 7046 9365 7098
rect 9417 7046 10856 7098
rect 1104 7024 10856 7046
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 9766 6984 9772 6996
rect 3660 6956 9772 6984
rect 3660 6944 3666 6956
rect 9766 6944 9772 6956
rect 9824 6944 9830 6996
rect 2133 6851 2191 6857
rect 2133 6817 2145 6851
rect 2179 6848 2191 6851
rect 3050 6848 3056 6860
rect 2179 6820 3056 6848
rect 2179 6817 2191 6820
rect 2133 6811 2191 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 2866 6740 2872 6792
rect 2924 6780 2930 6792
rect 2961 6783 3019 6789
rect 2961 6780 2973 6783
rect 2924 6752 2973 6780
rect 2924 6740 2930 6752
rect 2961 6749 2973 6752
rect 3007 6749 3019 6783
rect 3786 6780 3792 6792
rect 3747 6752 3792 6780
rect 2961 6743 3019 6749
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 1854 6712 1860 6724
rect 1815 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 6454 6712 6460 6724
rect 2792 6684 6460 6712
rect 2792 6653 2820 6684
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 2777 6647 2835 6653
rect 2777 6613 2789 6647
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 3050 6644 3056 6656
rect 2924 6616 3056 6644
rect 2924 6604 2930 6616
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 10042 6644 10048 6656
rect 10003 6616 10048 6644
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 1104 6554 10856 6576
rect 1104 6502 4213 6554
rect 4265 6502 4277 6554
rect 4329 6502 4341 6554
rect 4393 6502 4405 6554
rect 4457 6502 4469 6554
rect 4521 6502 7477 6554
rect 7529 6502 7541 6554
rect 7593 6502 7605 6554
rect 7657 6502 7669 6554
rect 7721 6502 7733 6554
rect 7785 6502 10856 6554
rect 1104 6480 10856 6502
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 4062 6440 4068 6452
rect 3283 6412 4068 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1964 6236 1992 6267
rect 2038 6264 2044 6316
rect 2096 6304 2102 6316
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 2096 6276 2605 6304
rect 2096 6264 2102 6276
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 2593 6267 2651 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3878 6236 3884 6248
rect 1964 6208 3884 6236
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6168 2835 6171
rect 9858 6168 9864 6180
rect 2823 6140 9864 6168
rect 2823 6137 2835 6140
rect 2777 6131 2835 6137
rect 9858 6128 9864 6140
rect 9916 6128 9922 6180
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 4798 6100 4804 6112
rect 2179 6072 4804 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 1104 6010 10856 6032
rect 1104 5958 2582 6010
rect 2634 5958 2646 6010
rect 2698 5958 2710 6010
rect 2762 5958 2774 6010
rect 2826 5958 2838 6010
rect 2890 5958 5845 6010
rect 5897 5958 5909 6010
rect 5961 5958 5973 6010
rect 6025 5958 6037 6010
rect 6089 5958 6101 6010
rect 6153 5958 9109 6010
rect 9161 5958 9173 6010
rect 9225 5958 9237 6010
rect 9289 5958 9301 6010
rect 9353 5958 9365 6010
rect 9417 5958 10856 6010
rect 1104 5936 10856 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 2958 5896 2964 5908
rect 2823 5868 2964 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3789 5899 3847 5905
rect 3789 5896 3801 5899
rect 3384 5868 3801 5896
rect 3384 5856 3390 5868
rect 3789 5865 3801 5868
rect 3835 5865 3847 5899
rect 3789 5859 3847 5865
rect 1489 5831 1547 5837
rect 1489 5797 1501 5831
rect 1535 5828 1547 5831
rect 6822 5828 6828 5840
rect 1535 5800 6828 5828
rect 1535 5797 1547 5800
rect 1489 5791 1547 5797
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 9674 5788 9680 5840
rect 9732 5788 9738 5840
rect 3050 5760 3056 5772
rect 2148 5732 3056 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2038 5692 2044 5704
rect 1719 5664 2044 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 2148 5701 2176 5732
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 9692 5760 9720 5788
rect 6886 5732 9720 5760
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2958 5692 2964 5704
rect 2919 5664 2964 5692
rect 2133 5655 2191 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 6886 5624 6914 5732
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 9861 5695 9919 5701
rect 9861 5692 9873 5695
rect 9732 5664 9873 5692
rect 9732 5652 9738 5664
rect 9861 5661 9873 5664
rect 9907 5661 9919 5695
rect 9861 5655 9919 5661
rect 2332 5596 6914 5624
rect 2332 5565 2360 5596
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5525 2375 5559
rect 10042 5556 10048 5568
rect 10003 5528 10048 5556
rect 2317 5519 2375 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 1104 5466 10856 5488
rect 1104 5414 4213 5466
rect 4265 5414 4277 5466
rect 4329 5414 4341 5466
rect 4393 5414 4405 5466
rect 4457 5414 4469 5466
rect 4521 5414 7477 5466
rect 7529 5414 7541 5466
rect 7593 5414 7605 5466
rect 7657 5414 7669 5466
rect 7721 5414 7733 5466
rect 7785 5414 10856 5466
rect 1104 5392 10856 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 3510 5352 3516 5364
rect 1995 5324 3516 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 3510 5312 3516 5324
rect 3568 5312 3574 5364
rect 1210 5244 1216 5296
rect 1268 5284 1274 5296
rect 1268 5256 3004 5284
rect 1268 5244 1274 5256
rect 2976 5225 3004 5256
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 2041 5179 2099 5185
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 3145 5219 3203 5225
rect 3145 5185 3157 5219
rect 3191 5216 3203 5219
rect 3234 5216 3240 5228
rect 3191 5188 3240 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 2056 5148 2084 5179
rect 3234 5176 3240 5188
rect 3292 5216 3298 5228
rect 3510 5216 3516 5228
rect 3292 5188 3516 5216
rect 3292 5176 3298 5188
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5216 9919 5219
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 9907 5188 11161 5216
rect 9907 5185 9919 5188
rect 9861 5179 9919 5185
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 3326 5148 3332 5160
rect 2056 5120 3332 5148
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3145 5015 3203 5021
rect 3145 4981 3157 5015
rect 3191 5012 3203 5015
rect 6362 5012 6368 5024
rect 3191 4984 6368 5012
rect 3191 4981 3203 4984
rect 3145 4975 3203 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 10042 5012 10048 5024
rect 10003 4984 10048 5012
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 1104 4922 10856 4944
rect 1104 4870 2582 4922
rect 2634 4870 2646 4922
rect 2698 4870 2710 4922
rect 2762 4870 2774 4922
rect 2826 4870 2838 4922
rect 2890 4870 5845 4922
rect 5897 4870 5909 4922
rect 5961 4870 5973 4922
rect 6025 4870 6037 4922
rect 6089 4870 6101 4922
rect 6153 4870 9109 4922
rect 9161 4870 9173 4922
rect 9225 4870 9237 4922
rect 9289 4870 9301 4922
rect 9353 4870 9365 4922
rect 9417 4870 10856 4922
rect 1104 4848 10856 4870
rect 3142 4768 3148 4820
rect 3200 4808 3206 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3200 4780 3801 4808
rect 3200 4768 3206 4780
rect 3789 4777 3801 4780
rect 3835 4777 3847 4811
rect 3789 4771 3847 4777
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 6270 4740 6276 4752
rect 1627 4712 6276 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1578 4604 1584 4616
rect 1443 4576 1584 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1578 4564 1584 4576
rect 1636 4604 1642 4616
rect 2409 4607 2467 4613
rect 2409 4604 2421 4607
rect 1636 4576 2421 4604
rect 1636 4564 1642 4576
rect 2409 4573 2421 4576
rect 2455 4573 2467 4607
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 2409 4567 2467 4573
rect 2516 4576 3065 4604
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 2516 4536 2544 4576
rect 3053 4573 3065 4576
rect 3099 4573 3111 4607
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 3053 4567 3111 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9824 4576 9873 4604
rect 9824 4564 9830 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 9674 4536 9680 4548
rect 1728 4508 2544 4536
rect 2608 4508 9680 4536
rect 1728 4496 1734 4508
rect 2608 4477 2636 4508
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4437 2651 4471
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 2593 4431 2651 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 10042 4468 10048 4480
rect 10003 4440 10048 4468
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 1104 4378 10856 4400
rect 1104 4326 4213 4378
rect 4265 4326 4277 4378
rect 4329 4326 4341 4378
rect 4393 4326 4405 4378
rect 4457 4326 4469 4378
rect 4521 4326 7477 4378
rect 7529 4326 7541 4378
rect 7593 4326 7605 4378
rect 7657 4326 7669 4378
rect 7721 4326 7733 4378
rect 7785 4326 10856 4378
rect 1104 4304 10856 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 9766 4264 9772 4276
rect 3292 4236 9772 4264
rect 3292 4224 3298 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 1210 4088 1216 4140
rect 1268 4128 1274 4140
rect 1857 4131 1915 4137
rect 1857 4128 1869 4131
rect 1268 4100 1869 4128
rect 1268 4088 1274 4100
rect 1857 4097 1869 4100
rect 1903 4097 1915 4131
rect 1857 4091 1915 4097
rect 2133 4131 2191 4137
rect 2133 4097 2145 4131
rect 2179 4128 2191 4131
rect 2222 4128 2228 4140
rect 2179 4100 2228 4128
rect 2179 4097 2191 4100
rect 2133 4091 2191 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2556 4100 2605 4128
rect 2556 4088 2562 4100
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 2915 4100 3341 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3510 4128 3516 4140
rect 3471 4100 3516 4128
rect 3329 4091 3387 4097
rect 3344 4060 3372 4091
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3602 4088 3608 4140
rect 3660 4128 3666 4140
rect 4157 4131 4215 4137
rect 4157 4128 4169 4131
rect 3660 4100 4169 4128
rect 3660 4088 3666 4100
rect 4157 4097 4169 4100
rect 4203 4097 4215 4131
rect 4157 4091 4215 4097
rect 5534 4060 5540 4072
rect 3344 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 9858 3992 9864 4004
rect 3559 3964 9864 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 3050 3884 3056 3936
rect 3108 3924 3114 3936
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3108 3896 3985 3924
rect 3108 3884 3114 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 3973 3887 4031 3893
rect 1104 3834 10856 3856
rect 1104 3782 2582 3834
rect 2634 3782 2646 3834
rect 2698 3782 2710 3834
rect 2762 3782 2774 3834
rect 2826 3782 2838 3834
rect 2890 3782 5845 3834
rect 5897 3782 5909 3834
rect 5961 3782 5973 3834
rect 6025 3782 6037 3834
rect 6089 3782 6101 3834
rect 6153 3782 9109 3834
rect 9161 3782 9173 3834
rect 9225 3782 9237 3834
rect 9289 3782 9301 3834
rect 9353 3782 9365 3834
rect 9417 3782 10856 3834
rect 1104 3760 10856 3782
rect 2225 3723 2283 3729
rect 2225 3689 2237 3723
rect 2271 3720 2283 3723
rect 2314 3720 2320 3732
rect 2271 3692 2320 3720
rect 2271 3689 2283 3692
rect 2225 3683 2283 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 1489 3655 1547 3661
rect 1489 3621 1501 3655
rect 1535 3652 1547 3655
rect 8110 3652 8116 3664
rect 1535 3624 8116 3652
rect 1535 3621 1547 3624
rect 1489 3615 1547 3621
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 1670 3516 1676 3528
rect 1631 3488 1676 3516
rect 1670 3476 1676 3488
rect 1728 3476 1734 3528
rect 2317 3519 2375 3525
rect 2317 3485 2329 3519
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 2332 3448 2360 3479
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 2961 3519 3019 3525
rect 2961 3516 2973 3519
rect 2464 3488 2973 3516
rect 2464 3476 2470 3488
rect 2961 3485 2973 3488
rect 3007 3485 3019 3519
rect 2961 3479 3019 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3510 3516 3516 3528
rect 3191 3488 3516 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 6886 3488 9873 3516
rect 3786 3448 3792 3460
rect 2332 3420 3792 3448
rect 3786 3408 3792 3420
rect 3844 3408 3850 3460
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 6886 3380 6914 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10042 3380 10048 3392
rect 3099 3352 6914 3380
rect 10003 3352 10048 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 1104 3290 10856 3312
rect 1104 3238 4213 3290
rect 4265 3238 4277 3290
rect 4329 3238 4341 3290
rect 4393 3238 4405 3290
rect 4457 3238 4469 3290
rect 4521 3238 7477 3290
rect 7529 3238 7541 3290
rect 7593 3238 7605 3290
rect 7657 3238 7669 3290
rect 7721 3238 7733 3290
rect 7785 3238 10856 3290
rect 1104 3216 10856 3238
rect 2222 3136 2228 3188
rect 2280 3176 2286 3188
rect 3973 3179 4031 3185
rect 3973 3176 3985 3179
rect 2280 3148 3985 3176
rect 2280 3136 2286 3148
rect 3973 3145 3985 3148
rect 4019 3145 4031 3179
rect 3973 3139 4031 3145
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2130 3040 2136 3052
rect 1719 3012 2136 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2866 3040 2872 3052
rect 2827 3012 2872 3040
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 3660 3012 4169 3040
rect 3660 3000 3666 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 6362 3000 6368 3052
rect 6420 3040 6426 3052
rect 9125 3043 9183 3049
rect 9125 3040 9137 3043
rect 6420 3012 9137 3040
rect 6420 3000 6426 3012
rect 9125 3009 9137 3012
rect 9171 3009 9183 3043
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9125 3003 9183 3009
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 2038 2864 2044 2916
rect 2096 2904 2102 2916
rect 2685 2907 2743 2913
rect 2685 2904 2697 2907
rect 2096 2876 2697 2904
rect 2096 2864 2102 2876
rect 2685 2873 2697 2876
rect 2731 2873 2743 2907
rect 3326 2904 3332 2916
rect 3287 2876 3332 2904
rect 2685 2867 2743 2873
rect 3326 2864 3332 2876
rect 3384 2864 3390 2916
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 9490 2836 9496 2848
rect 9355 2808 9496 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 1104 2746 10856 2768
rect 1104 2694 2582 2746
rect 2634 2694 2646 2746
rect 2698 2694 2710 2746
rect 2762 2694 2774 2746
rect 2826 2694 2838 2746
rect 2890 2694 5845 2746
rect 5897 2694 5909 2746
rect 5961 2694 5973 2746
rect 6025 2694 6037 2746
rect 6089 2694 6101 2746
rect 6153 2694 9109 2746
rect 9161 2694 9173 2746
rect 9225 2694 9237 2746
rect 9289 2694 9301 2746
rect 9353 2694 9365 2746
rect 9417 2694 10856 2746
rect 1104 2672 10856 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 1670 2592 1676 2644
rect 1728 2632 1734 2644
rect 2225 2635 2283 2641
rect 2225 2632 2237 2635
rect 1728 2604 2237 2632
rect 1728 2592 1734 2604
rect 2225 2601 2237 2604
rect 2271 2601 2283 2635
rect 2225 2595 2283 2601
rect 2498 2592 2504 2644
rect 2556 2632 2562 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2556 2604 2697 2632
rect 2556 2592 2562 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 2685 2595 2743 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 3936 2604 4445 2632
rect 3936 2592 3942 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2428 2099 2431
rect 2774 2428 2780 2440
rect 2087 2400 2780 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 2774 2388 2780 2400
rect 2832 2388 2838 2440
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 3970 2428 3976 2440
rect 2924 2400 2969 2428
rect 3931 2400 3976 2428
rect 2924 2388 2930 2400
rect 3970 2388 3976 2400
rect 4028 2388 4034 2440
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9824 2400 9873 2428
rect 9824 2388 9830 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 10042 2292 10048 2304
rect 10003 2264 10048 2292
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 1104 2202 10856 2224
rect 1104 2150 4213 2202
rect 4265 2150 4277 2202
rect 4329 2150 4341 2202
rect 4393 2150 4405 2202
rect 4457 2150 4469 2202
rect 4521 2150 7477 2202
rect 7529 2150 7541 2202
rect 7593 2150 7605 2202
rect 7657 2150 7669 2202
rect 7721 2150 7733 2202
rect 7785 2150 10856 2202
rect 1104 2128 10856 2150
rect 2774 484 2780 536
rect 2832 524 2838 536
rect 4614 524 4620 536
rect 2832 496 4620 524
rect 2832 484 2838 496
rect 4614 484 4620 496
rect 4672 484 4678 536
<< via1 >>
rect 10968 77979 11020 77988
rect 10968 77945 10977 77979
rect 10977 77945 11011 77979
rect 11011 77945 11020 77979
rect 10968 77936 11020 77945
rect 2582 77766 2634 77818
rect 2646 77766 2698 77818
rect 2710 77766 2762 77818
rect 2774 77766 2826 77818
rect 2838 77766 2890 77818
rect 5845 77766 5897 77818
rect 5909 77766 5961 77818
rect 5973 77766 6025 77818
rect 6037 77766 6089 77818
rect 6101 77766 6153 77818
rect 9109 77766 9161 77818
rect 9173 77766 9225 77818
rect 9237 77766 9289 77818
rect 9301 77766 9353 77818
rect 9365 77766 9417 77818
rect 3240 77596 3292 77648
rect 4712 77596 4764 77648
rect 3056 77528 3108 77580
rect 2504 77503 2556 77512
rect 2504 77469 2513 77503
rect 2513 77469 2547 77503
rect 2547 77469 2556 77503
rect 2504 77460 2556 77469
rect 3976 77503 4028 77512
rect 3976 77469 3985 77503
rect 3985 77469 4019 77503
rect 4019 77469 4028 77503
rect 3976 77460 4028 77469
rect 4068 77460 4120 77512
rect 9404 77503 9456 77512
rect 9404 77469 9413 77503
rect 9413 77469 9447 77503
rect 9447 77469 9456 77503
rect 9404 77460 9456 77469
rect 10140 77503 10192 77512
rect 10140 77469 10149 77503
rect 10149 77469 10183 77503
rect 10183 77469 10192 77503
rect 10140 77460 10192 77469
rect 1124 77392 1176 77444
rect 2964 77392 3016 77444
rect 3056 77324 3108 77376
rect 4620 77324 4672 77376
rect 5080 77367 5132 77376
rect 5080 77333 5089 77367
rect 5089 77333 5123 77367
rect 5123 77333 5132 77367
rect 5080 77324 5132 77333
rect 4213 77222 4265 77274
rect 4277 77222 4329 77274
rect 4341 77222 4393 77274
rect 4405 77222 4457 77274
rect 4469 77222 4521 77274
rect 7477 77222 7529 77274
rect 7541 77222 7593 77274
rect 7605 77222 7657 77274
rect 7669 77222 7721 77274
rect 7733 77222 7785 77274
rect 1400 77027 1452 77036
rect 1400 76993 1409 77027
rect 1409 76993 1443 77027
rect 1443 76993 1452 77027
rect 1400 76984 1452 76993
rect 2044 77027 2096 77036
rect 2044 76993 2053 77027
rect 2053 76993 2087 77027
rect 2087 76993 2096 77027
rect 2044 76984 2096 76993
rect 2780 76984 2832 77036
rect 3332 77027 3384 77036
rect 3332 76993 3341 77027
rect 3341 76993 3375 77027
rect 3375 76993 3384 77027
rect 3332 76984 3384 76993
rect 4160 77027 4212 77036
rect 4160 76993 4169 77027
rect 4169 76993 4203 77027
rect 4203 76993 4212 77027
rect 4160 76984 4212 76993
rect 10140 77027 10192 77036
rect 10140 76993 10149 77027
rect 10149 76993 10183 77027
rect 10183 76993 10192 77027
rect 10140 76984 10192 76993
rect 3424 76848 3476 76900
rect 1584 76823 1636 76832
rect 1584 76789 1593 76823
rect 1593 76789 1627 76823
rect 1627 76789 1636 76823
rect 1584 76780 1636 76789
rect 2228 76823 2280 76832
rect 2228 76789 2237 76823
rect 2237 76789 2271 76823
rect 2271 76789 2280 76823
rect 2228 76780 2280 76789
rect 3516 76823 3568 76832
rect 3516 76789 3525 76823
rect 3525 76789 3559 76823
rect 3559 76789 3568 76823
rect 3516 76780 3568 76789
rect 3976 76823 4028 76832
rect 3976 76789 3985 76823
rect 3985 76789 4019 76823
rect 4019 76789 4028 76823
rect 3976 76780 4028 76789
rect 9864 76780 9916 76832
rect 2582 76678 2634 76730
rect 2646 76678 2698 76730
rect 2710 76678 2762 76730
rect 2774 76678 2826 76730
rect 2838 76678 2890 76730
rect 5845 76678 5897 76730
rect 5909 76678 5961 76730
rect 5973 76678 6025 76730
rect 6037 76678 6089 76730
rect 6101 76678 6153 76730
rect 9109 76678 9161 76730
rect 9173 76678 9225 76730
rect 9237 76678 9289 76730
rect 9301 76678 9353 76730
rect 9365 76678 9417 76730
rect 1860 76576 1912 76628
rect 5080 76576 5132 76628
rect 1216 76508 1268 76560
rect 2780 76508 2832 76560
rect 3884 76508 3936 76560
rect 1676 76415 1728 76424
rect 1676 76381 1685 76415
rect 1685 76381 1719 76415
rect 1719 76381 1728 76415
rect 1676 76372 1728 76381
rect 3976 76440 4028 76492
rect 2136 76415 2188 76424
rect 2136 76381 2139 76415
rect 2139 76381 2188 76415
rect 2136 76372 2188 76381
rect 2780 76372 2832 76424
rect 2964 76415 3016 76424
rect 2964 76381 2973 76415
rect 2973 76381 3007 76415
rect 3007 76381 3016 76415
rect 2964 76372 3016 76381
rect 3148 76236 3200 76288
rect 4213 76134 4265 76186
rect 4277 76134 4329 76186
rect 4341 76134 4393 76186
rect 4405 76134 4457 76186
rect 4469 76134 4521 76186
rect 7477 76134 7529 76186
rect 7541 76134 7593 76186
rect 7605 76134 7657 76186
rect 7669 76134 7721 76186
rect 7733 76134 7785 76186
rect 1860 76007 1912 76016
rect 1860 75973 1869 76007
rect 1869 75973 1903 76007
rect 1903 75973 1912 76007
rect 1860 75964 1912 75973
rect 1676 75939 1728 75948
rect 1676 75905 1685 75939
rect 1685 75905 1719 75939
rect 1719 75905 1728 75939
rect 1676 75896 1728 75905
rect 2136 75939 2188 75948
rect 2136 75905 2139 75939
rect 2139 75905 2188 75939
rect 2136 75896 2188 75905
rect 4712 76032 4764 76084
rect 3608 75896 3660 75948
rect 6368 75896 6420 75948
rect 10232 75828 10284 75880
rect 1768 75692 1820 75744
rect 9956 75735 10008 75744
rect 9956 75701 9965 75735
rect 9965 75701 9999 75735
rect 9999 75701 10008 75735
rect 9956 75692 10008 75701
rect 2582 75590 2634 75642
rect 2646 75590 2698 75642
rect 2710 75590 2762 75642
rect 2774 75590 2826 75642
rect 2838 75590 2890 75642
rect 5845 75590 5897 75642
rect 5909 75590 5961 75642
rect 5973 75590 6025 75642
rect 6037 75590 6089 75642
rect 6101 75590 6153 75642
rect 9109 75590 9161 75642
rect 9173 75590 9225 75642
rect 9237 75590 9289 75642
rect 9301 75590 9353 75642
rect 9365 75590 9417 75642
rect 388 75420 440 75472
rect 1308 75284 1360 75336
rect 2596 75327 2648 75336
rect 2596 75293 2600 75327
rect 2600 75293 2634 75327
rect 2634 75293 2648 75327
rect 2596 75284 2648 75293
rect 2964 75327 3016 75336
rect 2964 75293 2973 75327
rect 2973 75293 3007 75327
rect 3007 75293 3016 75327
rect 3976 75327 4028 75336
rect 2964 75284 3016 75293
rect 3976 75293 3985 75327
rect 3985 75293 4019 75327
rect 4019 75293 4028 75327
rect 3976 75284 4028 75293
rect 10140 75327 10192 75336
rect 10140 75293 10149 75327
rect 10149 75293 10183 75327
rect 10183 75293 10192 75327
rect 10140 75284 10192 75293
rect 1860 75148 1912 75200
rect 3056 75148 3108 75200
rect 3792 75191 3844 75200
rect 3792 75157 3801 75191
rect 3801 75157 3835 75191
rect 3835 75157 3844 75191
rect 3792 75148 3844 75157
rect 4213 75046 4265 75098
rect 4277 75046 4329 75098
rect 4341 75046 4393 75098
rect 4405 75046 4457 75098
rect 4469 75046 4521 75098
rect 7477 75046 7529 75098
rect 7541 75046 7593 75098
rect 7605 75046 7657 75098
rect 7669 75046 7721 75098
rect 7733 75046 7785 75098
rect 2872 74944 2924 74996
rect 4620 74944 4672 74996
rect 1400 74851 1452 74860
rect 1400 74817 1409 74851
rect 1409 74817 1443 74851
rect 1443 74817 1452 74851
rect 1400 74808 1452 74817
rect 2596 74851 2648 74860
rect 2596 74817 2600 74851
rect 2600 74817 2634 74851
rect 2634 74817 2648 74851
rect 2596 74808 2648 74817
rect 2872 74808 2924 74860
rect 2964 74851 3016 74860
rect 2964 74817 2973 74851
rect 2973 74817 3007 74851
rect 3007 74817 3016 74851
rect 2964 74808 3016 74817
rect 3332 74808 3384 74860
rect 3516 74876 3568 74928
rect 9864 74876 9916 74928
rect 3884 74851 3936 74860
rect 3884 74817 3887 74851
rect 3887 74817 3936 74851
rect 3884 74808 3936 74817
rect 9956 74740 10008 74792
rect 1952 74604 2004 74656
rect 4620 74672 4672 74724
rect 8300 74604 8352 74656
rect 2582 74502 2634 74554
rect 2646 74502 2698 74554
rect 2710 74502 2762 74554
rect 2774 74502 2826 74554
rect 2838 74502 2890 74554
rect 5845 74502 5897 74554
rect 5909 74502 5961 74554
rect 5973 74502 6025 74554
rect 6037 74502 6089 74554
rect 6101 74502 6153 74554
rect 9109 74502 9161 74554
rect 9173 74502 9225 74554
rect 9237 74502 9289 74554
rect 9301 74502 9353 74554
rect 9365 74502 9417 74554
rect 1584 74239 1636 74248
rect 1584 74205 1593 74239
rect 1593 74205 1627 74239
rect 1627 74205 1636 74239
rect 1584 74196 1636 74205
rect 4896 74332 4948 74384
rect 1492 74128 1544 74180
rect 2504 74196 2556 74248
rect 2780 74196 2832 74248
rect 3332 74196 3384 74248
rect 10140 74239 10192 74248
rect 10140 74205 10149 74239
rect 10149 74205 10183 74239
rect 10183 74205 10192 74239
rect 10140 74196 10192 74205
rect 2136 74060 2188 74112
rect 3240 74060 3292 74112
rect 9772 74060 9824 74112
rect 4213 73958 4265 74010
rect 4277 73958 4329 74010
rect 4341 73958 4393 74010
rect 4405 73958 4457 74010
rect 4469 73958 4521 74010
rect 7477 73958 7529 74010
rect 7541 73958 7593 74010
rect 7605 73958 7657 74010
rect 7669 73958 7721 74010
rect 7733 73958 7785 74010
rect 3148 73788 3200 73840
rect 1492 73720 1544 73772
rect 2136 73720 2188 73772
rect 2964 73720 3016 73772
rect 10140 73763 10192 73772
rect 10140 73729 10149 73763
rect 10149 73729 10183 73763
rect 10183 73729 10192 73763
rect 10140 73720 10192 73729
rect 9956 73652 10008 73704
rect 5540 73584 5592 73636
rect 2320 73516 2372 73568
rect 2582 73414 2634 73466
rect 2646 73414 2698 73466
rect 2710 73414 2762 73466
rect 2774 73414 2826 73466
rect 2838 73414 2890 73466
rect 5845 73414 5897 73466
rect 5909 73414 5961 73466
rect 5973 73414 6025 73466
rect 6037 73414 6089 73466
rect 6101 73414 6153 73466
rect 9109 73414 9161 73466
rect 9173 73414 9225 73466
rect 9237 73414 9289 73466
rect 9301 73414 9353 73466
rect 9365 73414 9417 73466
rect 1400 73151 1452 73160
rect 1400 73117 1409 73151
rect 1409 73117 1443 73151
rect 1443 73117 1452 73151
rect 1400 73108 1452 73117
rect 2228 73151 2280 73160
rect 2228 73117 2237 73151
rect 2237 73117 2271 73151
rect 2271 73117 2280 73151
rect 2228 73108 2280 73117
rect 10140 73151 10192 73160
rect 10140 73117 10149 73151
rect 10149 73117 10183 73151
rect 10183 73117 10192 73151
rect 10140 73108 10192 73117
rect 1676 72972 1728 73024
rect 2044 73015 2096 73024
rect 2044 72981 2053 73015
rect 2053 72981 2087 73015
rect 2087 72981 2096 73015
rect 2044 72972 2096 72981
rect 4213 72870 4265 72922
rect 4277 72870 4329 72922
rect 4341 72870 4393 72922
rect 4405 72870 4457 72922
rect 4469 72870 4521 72922
rect 7477 72870 7529 72922
rect 7541 72870 7593 72922
rect 7605 72870 7657 72922
rect 7669 72870 7721 72922
rect 7733 72870 7785 72922
rect 1308 72632 1360 72684
rect 2228 72428 2280 72480
rect 2582 72326 2634 72378
rect 2646 72326 2698 72378
rect 2710 72326 2762 72378
rect 2774 72326 2826 72378
rect 2838 72326 2890 72378
rect 5845 72326 5897 72378
rect 5909 72326 5961 72378
rect 5973 72326 6025 72378
rect 6037 72326 6089 72378
rect 6101 72326 6153 72378
rect 9109 72326 9161 72378
rect 9173 72326 9225 72378
rect 9237 72326 9289 72378
rect 9301 72326 9353 72378
rect 9365 72326 9417 72378
rect 1400 72224 1452 72276
rect 2136 72224 2188 72276
rect 9956 72267 10008 72276
rect 9956 72233 9965 72267
rect 9965 72233 9999 72267
rect 9999 72233 10008 72267
rect 9956 72224 10008 72233
rect 1400 72063 1452 72072
rect 1400 72029 1409 72063
rect 1409 72029 1443 72063
rect 1443 72029 1452 72063
rect 1400 72020 1452 72029
rect 3792 72088 3844 72140
rect 1768 72020 1820 72072
rect 3240 72020 3292 72072
rect 10140 72063 10192 72072
rect 10140 72029 10149 72063
rect 10149 72029 10183 72063
rect 10183 72029 10192 72063
rect 10140 72020 10192 72029
rect 9864 71952 9916 72004
rect 1492 71884 1544 71936
rect 1768 71884 1820 71936
rect 4213 71782 4265 71834
rect 4277 71782 4329 71834
rect 4341 71782 4393 71834
rect 4405 71782 4457 71834
rect 4469 71782 4521 71834
rect 7477 71782 7529 71834
rect 7541 71782 7593 71834
rect 7605 71782 7657 71834
rect 7669 71782 7721 71834
rect 7733 71782 7785 71834
rect 9772 71680 9824 71732
rect 10140 71587 10192 71596
rect 10140 71553 10149 71587
rect 10149 71553 10183 71587
rect 10183 71553 10192 71587
rect 10140 71544 10192 71553
rect 1400 71519 1452 71528
rect 1400 71485 1409 71519
rect 1409 71485 1443 71519
rect 1443 71485 1452 71519
rect 1400 71476 1452 71485
rect 1768 71476 1820 71528
rect 2582 71238 2634 71290
rect 2646 71238 2698 71290
rect 2710 71238 2762 71290
rect 2774 71238 2826 71290
rect 2838 71238 2890 71290
rect 5845 71238 5897 71290
rect 5909 71238 5961 71290
rect 5973 71238 6025 71290
rect 6037 71238 6089 71290
rect 6101 71238 6153 71290
rect 9109 71238 9161 71290
rect 9173 71238 9225 71290
rect 9237 71238 9289 71290
rect 9301 71238 9353 71290
rect 9365 71238 9417 71290
rect 1308 71000 1360 71052
rect 2504 70932 2556 70984
rect 2780 70932 2832 70984
rect 4068 70796 4120 70848
rect 4213 70694 4265 70746
rect 4277 70694 4329 70746
rect 4341 70694 4393 70746
rect 4405 70694 4457 70746
rect 4469 70694 4521 70746
rect 7477 70694 7529 70746
rect 7541 70694 7593 70746
rect 7605 70694 7657 70746
rect 7669 70694 7721 70746
rect 7733 70694 7785 70746
rect 2688 70592 2740 70644
rect 2872 70592 2924 70644
rect 3424 70592 3476 70644
rect 9864 70592 9916 70644
rect 940 70320 992 70372
rect 1768 70320 1820 70372
rect 1584 70295 1636 70304
rect 1584 70261 1593 70295
rect 1593 70261 1627 70295
rect 1627 70261 1636 70295
rect 1584 70252 1636 70261
rect 2780 70456 2832 70508
rect 2964 70456 3016 70508
rect 3332 70456 3384 70508
rect 3516 70499 3568 70508
rect 3516 70465 3525 70499
rect 3525 70465 3559 70499
rect 3559 70465 3568 70499
rect 3516 70456 3568 70465
rect 10140 70499 10192 70508
rect 10140 70465 10149 70499
rect 10149 70465 10183 70499
rect 10183 70465 10192 70499
rect 10140 70456 10192 70465
rect 7012 70388 7064 70440
rect 2780 70320 2832 70372
rect 3148 70320 3200 70372
rect 3056 70252 3108 70304
rect 3608 70252 3660 70304
rect 2582 70150 2634 70202
rect 2646 70150 2698 70202
rect 2710 70150 2762 70202
rect 2774 70150 2826 70202
rect 2838 70150 2890 70202
rect 5845 70150 5897 70202
rect 5909 70150 5961 70202
rect 5973 70150 6025 70202
rect 6037 70150 6089 70202
rect 6101 70150 6153 70202
rect 9109 70150 9161 70202
rect 9173 70150 9225 70202
rect 9237 70150 9289 70202
rect 9301 70150 9353 70202
rect 9365 70150 9417 70202
rect 1308 69844 1360 69896
rect 2872 69912 2924 69964
rect 3056 69912 3108 69964
rect 2412 69776 2464 69828
rect 3240 69844 3292 69896
rect 3976 69887 4028 69896
rect 3976 69853 3985 69887
rect 3985 69853 4019 69887
rect 4019 69853 4028 69887
rect 3976 69844 4028 69853
rect 10140 69887 10192 69896
rect 10140 69853 10149 69887
rect 10149 69853 10183 69887
rect 10183 69853 10192 69887
rect 10140 69844 10192 69853
rect 3516 69708 3568 69760
rect 3700 69708 3752 69760
rect 9956 69751 10008 69760
rect 9956 69717 9965 69751
rect 9965 69717 9999 69751
rect 9999 69717 10008 69751
rect 9956 69708 10008 69717
rect 4213 69606 4265 69658
rect 4277 69606 4329 69658
rect 4341 69606 4393 69658
rect 4405 69606 4457 69658
rect 4469 69606 4521 69658
rect 7477 69606 7529 69658
rect 7541 69606 7593 69658
rect 7605 69606 7657 69658
rect 7669 69606 7721 69658
rect 7733 69606 7785 69658
rect 1584 69504 1636 69556
rect 3332 69504 3384 69556
rect 1768 69479 1820 69488
rect 1768 69445 1777 69479
rect 1777 69445 1811 69479
rect 1811 69445 1820 69479
rect 1768 69436 1820 69445
rect 1584 69368 1636 69420
rect 2136 69436 2188 69488
rect 5724 69436 5776 69488
rect 9956 69436 10008 69488
rect 2412 69368 2464 69420
rect 2964 69368 3016 69420
rect 3240 69368 3292 69420
rect 4160 69368 4212 69420
rect 10140 69411 10192 69420
rect 10140 69377 10149 69411
rect 10149 69377 10183 69411
rect 10183 69377 10192 69411
rect 10140 69368 10192 69377
rect 1768 69300 1820 69352
rect 3148 69300 3200 69352
rect 1400 69232 1452 69284
rect 1492 69207 1544 69216
rect 1492 69173 1501 69207
rect 1501 69173 1535 69207
rect 1535 69173 1544 69207
rect 1492 69164 1544 69173
rect 9956 69207 10008 69216
rect 9956 69173 9965 69207
rect 9965 69173 9999 69207
rect 9999 69173 10008 69207
rect 9956 69164 10008 69173
rect 2582 69062 2634 69114
rect 2646 69062 2698 69114
rect 2710 69062 2762 69114
rect 2774 69062 2826 69114
rect 2838 69062 2890 69114
rect 5845 69062 5897 69114
rect 5909 69062 5961 69114
rect 5973 69062 6025 69114
rect 6037 69062 6089 69114
rect 6101 69062 6153 69114
rect 9109 69062 9161 69114
rect 9173 69062 9225 69114
rect 9237 69062 9289 69114
rect 9301 69062 9353 69114
rect 9365 69062 9417 69114
rect 2964 68867 3016 68876
rect 2964 68833 2973 68867
rect 2973 68833 3007 68867
rect 3007 68833 3016 68867
rect 2964 68824 3016 68833
rect 1308 68756 1360 68808
rect 3976 68799 4028 68808
rect 2964 68688 3016 68740
rect 3976 68765 3985 68799
rect 3985 68765 4019 68799
rect 4019 68765 4028 68799
rect 3976 68756 4028 68765
rect 2136 68620 2188 68672
rect 3792 68663 3844 68672
rect 3792 68629 3801 68663
rect 3801 68629 3835 68663
rect 3835 68629 3844 68663
rect 3792 68620 3844 68629
rect 4213 68518 4265 68570
rect 4277 68518 4329 68570
rect 4341 68518 4393 68570
rect 4405 68518 4457 68570
rect 4469 68518 4521 68570
rect 7477 68518 7529 68570
rect 7541 68518 7593 68570
rect 7605 68518 7657 68570
rect 7669 68518 7721 68570
rect 7733 68518 7785 68570
rect 1860 68416 1912 68468
rect 1952 68391 2004 68400
rect 1952 68357 1961 68391
rect 1961 68357 1995 68391
rect 1995 68357 2004 68391
rect 1952 68348 2004 68357
rect 3240 68416 3292 68468
rect 1676 68280 1728 68332
rect 1492 68212 1544 68264
rect 9956 68348 10008 68400
rect 2412 68280 2464 68332
rect 3332 68323 3384 68332
rect 3332 68289 3335 68323
rect 3335 68289 3384 68323
rect 3332 68280 3384 68289
rect 3424 68280 3476 68332
rect 10140 68323 10192 68332
rect 10140 68289 10149 68323
rect 10149 68289 10183 68323
rect 10183 68289 10192 68323
rect 10140 68280 10192 68289
rect 7104 68212 7156 68264
rect 8484 68076 8536 68128
rect 2582 67974 2634 68026
rect 2646 67974 2698 68026
rect 2710 67974 2762 68026
rect 2774 67974 2826 68026
rect 2838 67974 2890 68026
rect 5845 67974 5897 68026
rect 5909 67974 5961 68026
rect 5973 67974 6025 68026
rect 6037 67974 6089 68026
rect 6101 67974 6153 68026
rect 9109 67974 9161 68026
rect 9173 67974 9225 68026
rect 9237 67974 9289 68026
rect 9301 67974 9353 68026
rect 9365 67974 9417 68026
rect 3792 67872 3844 67924
rect 1400 67804 1452 67856
rect 3148 67804 3200 67856
rect 3424 67804 3476 67856
rect 1400 67711 1452 67720
rect 1400 67677 1409 67711
rect 1409 67677 1443 67711
rect 1443 67677 1452 67711
rect 1400 67668 1452 67677
rect 1860 67668 1912 67720
rect 2964 67643 3016 67652
rect 2964 67609 2973 67643
rect 2973 67609 3007 67643
rect 3007 67609 3016 67643
rect 2964 67600 3016 67609
rect 3056 67600 3108 67652
rect 3884 67600 3936 67652
rect 9956 67575 10008 67584
rect 9956 67541 9965 67575
rect 9965 67541 9999 67575
rect 9999 67541 10008 67575
rect 9956 67532 10008 67541
rect 10140 67532 10192 67584
rect 4213 67430 4265 67482
rect 4277 67430 4329 67482
rect 4341 67430 4393 67482
rect 4405 67430 4457 67482
rect 4469 67430 4521 67482
rect 7477 67430 7529 67482
rect 7541 67430 7593 67482
rect 7605 67430 7657 67482
rect 7669 67430 7721 67482
rect 7733 67430 7785 67482
rect 3332 67328 3384 67380
rect 9956 67260 10008 67312
rect 1492 67192 1544 67244
rect 2320 67192 2372 67244
rect 1676 67124 1728 67176
rect 2964 67192 3016 67244
rect 3148 67192 3200 67244
rect 5356 67056 5408 67108
rect 2582 66886 2634 66938
rect 2646 66886 2698 66938
rect 2710 66886 2762 66938
rect 2774 66886 2826 66938
rect 2838 66886 2890 66938
rect 5845 66886 5897 66938
rect 5909 66886 5961 66938
rect 5973 66886 6025 66938
rect 6037 66886 6089 66938
rect 6101 66886 6153 66938
rect 9109 66886 9161 66938
rect 9173 66886 9225 66938
rect 9237 66886 9289 66938
rect 9301 66886 9353 66938
rect 9365 66886 9417 66938
rect 2320 66623 2372 66632
rect 2320 66589 2329 66623
rect 2329 66589 2363 66623
rect 2363 66589 2372 66623
rect 2320 66580 2372 66589
rect 2964 66623 3016 66632
rect 2964 66589 2973 66623
rect 2973 66589 3007 66623
rect 3007 66589 3016 66623
rect 2964 66580 3016 66589
rect 3332 66580 3384 66632
rect 3608 66580 3660 66632
rect 10140 66623 10192 66632
rect 10140 66589 10149 66623
rect 10149 66589 10183 66623
rect 10183 66589 10192 66623
rect 10140 66580 10192 66589
rect 6920 66512 6972 66564
rect 1492 66487 1544 66496
rect 1492 66453 1501 66487
rect 1501 66453 1535 66487
rect 1535 66453 1544 66487
rect 1492 66444 1544 66453
rect 2136 66487 2188 66496
rect 2136 66453 2145 66487
rect 2145 66453 2179 66487
rect 2179 66453 2188 66487
rect 2136 66444 2188 66453
rect 3608 66444 3660 66496
rect 9956 66487 10008 66496
rect 9956 66453 9965 66487
rect 9965 66453 9999 66487
rect 9999 66453 10008 66487
rect 9956 66444 10008 66453
rect 4213 66342 4265 66394
rect 4277 66342 4329 66394
rect 4341 66342 4393 66394
rect 4405 66342 4457 66394
rect 4469 66342 4521 66394
rect 7477 66342 7529 66394
rect 7541 66342 7593 66394
rect 7605 66342 7657 66394
rect 7669 66342 7721 66394
rect 7733 66342 7785 66394
rect 10140 66147 10192 66156
rect 10140 66113 10149 66147
rect 10149 66113 10183 66147
rect 10183 66113 10192 66147
rect 10140 66104 10192 66113
rect 1400 66079 1452 66088
rect 1400 66045 1409 66079
rect 1409 66045 1443 66079
rect 1443 66045 1452 66079
rect 1400 66036 1452 66045
rect 9864 65900 9916 65952
rect 2582 65798 2634 65850
rect 2646 65798 2698 65850
rect 2710 65798 2762 65850
rect 2774 65798 2826 65850
rect 2838 65798 2890 65850
rect 5845 65798 5897 65850
rect 5909 65798 5961 65850
rect 5973 65798 6025 65850
rect 6037 65798 6089 65850
rect 6101 65798 6153 65850
rect 9109 65798 9161 65850
rect 9173 65798 9225 65850
rect 9237 65798 9289 65850
rect 9301 65798 9353 65850
rect 9365 65798 9417 65850
rect 1032 65492 1084 65544
rect 480 65424 532 65476
rect 5632 65492 5684 65544
rect 10140 65535 10192 65544
rect 10140 65501 10149 65535
rect 10149 65501 10183 65535
rect 10183 65501 10192 65535
rect 10140 65492 10192 65501
rect 1492 65399 1544 65408
rect 1492 65365 1501 65399
rect 1501 65365 1535 65399
rect 1535 65365 1544 65399
rect 1492 65356 1544 65365
rect 2320 65399 2372 65408
rect 2320 65365 2329 65399
rect 2329 65365 2363 65399
rect 2363 65365 2372 65399
rect 2320 65356 2372 65365
rect 3056 65399 3108 65408
rect 3056 65365 3065 65399
rect 3065 65365 3099 65399
rect 3099 65365 3108 65399
rect 3056 65356 3108 65365
rect 9772 65356 9824 65408
rect 4213 65254 4265 65306
rect 4277 65254 4329 65306
rect 4341 65254 4393 65306
rect 4405 65254 4457 65306
rect 4469 65254 4521 65306
rect 7477 65254 7529 65306
rect 7541 65254 7593 65306
rect 7605 65254 7657 65306
rect 7669 65254 7721 65306
rect 7733 65254 7785 65306
rect 1952 65127 2004 65136
rect 1952 65093 1961 65127
rect 1961 65093 1995 65127
rect 1995 65093 2004 65127
rect 1952 65084 2004 65093
rect 9956 65084 10008 65136
rect 1676 65016 1728 65068
rect 1400 64948 1452 65000
rect 1952 64948 2004 65000
rect 3056 64948 3108 65000
rect 2582 64710 2634 64762
rect 2646 64710 2698 64762
rect 2710 64710 2762 64762
rect 2774 64710 2826 64762
rect 2838 64710 2890 64762
rect 5845 64710 5897 64762
rect 5909 64710 5961 64762
rect 5973 64710 6025 64762
rect 6037 64710 6089 64762
rect 6101 64710 6153 64762
rect 9109 64710 9161 64762
rect 9173 64710 9225 64762
rect 9237 64710 9289 64762
rect 9301 64710 9353 64762
rect 9365 64710 9417 64762
rect 1676 64540 1728 64592
rect 2412 64472 2464 64524
rect 10140 64447 10192 64456
rect 1400 64268 1452 64320
rect 10140 64413 10149 64447
rect 10149 64413 10183 64447
rect 10183 64413 10192 64447
rect 10140 64404 10192 64413
rect 3424 64336 3476 64388
rect 3792 64268 3844 64320
rect 4213 64166 4265 64218
rect 4277 64166 4329 64218
rect 4341 64166 4393 64218
rect 4405 64166 4457 64218
rect 4469 64166 4521 64218
rect 7477 64166 7529 64218
rect 7541 64166 7593 64218
rect 7605 64166 7657 64218
rect 7669 64166 7721 64218
rect 7733 64166 7785 64218
rect 9864 64064 9916 64116
rect 1952 63928 2004 63980
rect 1584 63860 1636 63912
rect 2412 63928 2464 63980
rect 5080 63928 5132 63980
rect 5172 63860 5224 63912
rect 10140 63903 10192 63912
rect 10140 63869 10149 63903
rect 10149 63869 10183 63903
rect 10183 63869 10192 63903
rect 10140 63860 10192 63869
rect 3884 63835 3936 63844
rect 3148 63767 3200 63776
rect 3148 63733 3157 63767
rect 3157 63733 3191 63767
rect 3191 63733 3200 63767
rect 3148 63724 3200 63733
rect 3884 63801 3893 63835
rect 3893 63801 3927 63835
rect 3927 63801 3936 63835
rect 3884 63792 3936 63801
rect 6276 63724 6328 63776
rect 2582 63622 2634 63674
rect 2646 63622 2698 63674
rect 2710 63622 2762 63674
rect 2774 63622 2826 63674
rect 2838 63622 2890 63674
rect 5845 63622 5897 63674
rect 5909 63622 5961 63674
rect 5973 63622 6025 63674
rect 6037 63622 6089 63674
rect 6101 63622 6153 63674
rect 9109 63622 9161 63674
rect 9173 63622 9225 63674
rect 9237 63622 9289 63674
rect 9301 63622 9353 63674
rect 9365 63622 9417 63674
rect 5448 63520 5500 63572
rect 8576 63452 8628 63504
rect 1676 63384 1728 63436
rect 2872 63384 2924 63436
rect 1952 63316 2004 63368
rect 2412 63316 2464 63368
rect 1676 63291 1728 63300
rect 1676 63257 1685 63291
rect 1685 63257 1719 63291
rect 1719 63257 1728 63291
rect 2872 63291 2924 63300
rect 1676 63248 1728 63257
rect 2872 63257 2881 63291
rect 2881 63257 2915 63291
rect 2915 63257 2924 63291
rect 2872 63248 2924 63257
rect 5724 63316 5776 63368
rect 3884 63248 3936 63300
rect 4068 63248 4120 63300
rect 9956 63248 10008 63300
rect 2320 63180 2372 63232
rect 3976 63223 4028 63232
rect 3976 63189 3985 63223
rect 3985 63189 4019 63223
rect 4019 63189 4028 63223
rect 3976 63180 4028 63189
rect 4213 63078 4265 63130
rect 4277 63078 4329 63130
rect 4341 63078 4393 63130
rect 4405 63078 4457 63130
rect 4469 63078 4521 63130
rect 7477 63078 7529 63130
rect 7541 63078 7593 63130
rect 7605 63078 7657 63130
rect 7669 63078 7721 63130
rect 7733 63078 7785 63130
rect 1676 62976 1728 63028
rect 9956 63019 10008 63028
rect 2320 62908 2372 62960
rect 9956 62985 9965 63019
rect 9965 62985 9999 63019
rect 9999 62985 10008 63019
rect 9956 62976 10008 62985
rect 1584 62840 1636 62892
rect 9772 62908 9824 62960
rect 940 62772 992 62824
rect 2320 62772 2372 62824
rect 1492 62679 1544 62688
rect 1492 62645 1501 62679
rect 1501 62645 1535 62679
rect 1535 62645 1544 62679
rect 1492 62636 1544 62645
rect 2228 62679 2280 62688
rect 2228 62645 2237 62679
rect 2237 62645 2271 62679
rect 2271 62645 2280 62679
rect 2228 62636 2280 62645
rect 4988 62840 5040 62892
rect 10140 62883 10192 62892
rect 10140 62849 10149 62883
rect 10149 62849 10183 62883
rect 10183 62849 10192 62883
rect 10140 62840 10192 62849
rect 3056 62772 3108 62824
rect 5448 62704 5500 62756
rect 3056 62636 3108 62688
rect 2582 62534 2634 62586
rect 2646 62534 2698 62586
rect 2710 62534 2762 62586
rect 2774 62534 2826 62586
rect 2838 62534 2890 62586
rect 5845 62534 5897 62586
rect 5909 62534 5961 62586
rect 5973 62534 6025 62586
rect 6037 62534 6089 62586
rect 6101 62534 6153 62586
rect 9109 62534 9161 62586
rect 9173 62534 9225 62586
rect 9237 62534 9289 62586
rect 9301 62534 9353 62586
rect 9365 62534 9417 62586
rect 664 62432 716 62484
rect 5448 62432 5500 62484
rect 1400 62364 1452 62416
rect 1768 62364 1820 62416
rect 9680 62296 9732 62348
rect 1768 62271 1820 62280
rect 1768 62237 1782 62271
rect 1782 62237 1816 62271
rect 1816 62237 1820 62271
rect 1768 62228 1820 62237
rect 2412 62228 2464 62280
rect 3884 62228 3936 62280
rect 10140 62271 10192 62280
rect 10140 62237 10149 62271
rect 10149 62237 10183 62271
rect 10183 62237 10192 62271
rect 10140 62228 10192 62237
rect 1952 62092 2004 62144
rect 3516 62160 3568 62212
rect 4213 61990 4265 62042
rect 4277 61990 4329 62042
rect 4341 61990 4393 62042
rect 4405 61990 4457 62042
rect 4469 61990 4521 62042
rect 7477 61990 7529 62042
rect 7541 61990 7593 62042
rect 7605 61990 7657 62042
rect 7669 61990 7721 62042
rect 7733 61990 7785 62042
rect 4068 61888 4120 61940
rect 2964 61820 3016 61872
rect 3148 61820 3200 61872
rect 1768 61795 1820 61804
rect 1768 61761 1782 61795
rect 1782 61761 1816 61795
rect 1816 61761 1820 61795
rect 1768 61752 1820 61761
rect 2044 61752 2096 61804
rect 10140 61795 10192 61804
rect 10140 61761 10149 61795
rect 10149 61761 10183 61795
rect 10183 61761 10192 61795
rect 10140 61752 10192 61761
rect 9772 61684 9824 61736
rect 3700 61616 3752 61668
rect 1952 61548 2004 61600
rect 2964 61548 3016 61600
rect 9956 61591 10008 61600
rect 9956 61557 9965 61591
rect 9965 61557 9999 61591
rect 9999 61557 10008 61591
rect 9956 61548 10008 61557
rect 2582 61446 2634 61498
rect 2646 61446 2698 61498
rect 2710 61446 2762 61498
rect 2774 61446 2826 61498
rect 2838 61446 2890 61498
rect 5845 61446 5897 61498
rect 5909 61446 5961 61498
rect 5973 61446 6025 61498
rect 6037 61446 6089 61498
rect 6101 61446 6153 61498
rect 9109 61446 9161 61498
rect 9173 61446 9225 61498
rect 9237 61446 9289 61498
rect 9301 61446 9353 61498
rect 9365 61446 9417 61498
rect 1768 61344 1820 61396
rect 2136 61344 2188 61396
rect 1952 61208 2004 61260
rect 1676 61183 1728 61192
rect 1676 61149 1680 61183
rect 1680 61149 1714 61183
rect 1714 61149 1728 61183
rect 1676 61140 1728 61149
rect 2228 61140 2280 61192
rect 3424 61140 3476 61192
rect 9864 61072 9916 61124
rect 2780 61004 2832 61056
rect 3976 61047 4028 61056
rect 3976 61013 3985 61047
rect 3985 61013 4019 61047
rect 4019 61013 4028 61047
rect 3976 61004 4028 61013
rect 4213 60902 4265 60954
rect 4277 60902 4329 60954
rect 4341 60902 4393 60954
rect 4405 60902 4457 60954
rect 4469 60902 4521 60954
rect 7477 60902 7529 60954
rect 7541 60902 7593 60954
rect 7605 60902 7657 60954
rect 7669 60902 7721 60954
rect 7733 60902 7785 60954
rect 1400 60800 1452 60852
rect 1860 60800 1912 60852
rect 2412 60800 2464 60852
rect 1584 60732 1636 60784
rect 3332 60800 3384 60852
rect 1308 60664 1360 60716
rect 1860 60664 1912 60716
rect 1492 60503 1544 60512
rect 1492 60469 1501 60503
rect 1501 60469 1535 60503
rect 1535 60469 1544 60503
rect 1492 60460 1544 60469
rect 9956 60732 10008 60784
rect 3608 60664 3660 60716
rect 10140 60707 10192 60716
rect 10140 60673 10149 60707
rect 10149 60673 10183 60707
rect 10183 60673 10192 60707
rect 10140 60664 10192 60673
rect 3332 60596 3384 60648
rect 9772 60528 9824 60580
rect 2320 60460 2372 60512
rect 3516 60460 3568 60512
rect 3608 60460 3660 60512
rect 2582 60358 2634 60410
rect 2646 60358 2698 60410
rect 2710 60358 2762 60410
rect 2774 60358 2826 60410
rect 2838 60358 2890 60410
rect 5845 60358 5897 60410
rect 5909 60358 5961 60410
rect 5973 60358 6025 60410
rect 6037 60358 6089 60410
rect 6101 60358 6153 60410
rect 9109 60358 9161 60410
rect 9173 60358 9225 60410
rect 9237 60358 9289 60410
rect 9301 60358 9353 60410
rect 9365 60358 9417 60410
rect 1860 60256 1912 60308
rect 3976 60256 4028 60308
rect 9680 60256 9732 60308
rect 1676 60188 1728 60240
rect 1308 59916 1360 59968
rect 1952 60052 2004 60104
rect 10140 60095 10192 60104
rect 10140 60061 10149 60095
rect 10149 60061 10183 60095
rect 10183 60061 10192 60095
rect 10140 60052 10192 60061
rect 2964 59984 3016 60036
rect 3148 59984 3200 60036
rect 2872 59916 2924 59968
rect 4213 59814 4265 59866
rect 4277 59814 4329 59866
rect 4341 59814 4393 59866
rect 4405 59814 4457 59866
rect 4469 59814 4521 59866
rect 7477 59814 7529 59866
rect 7541 59814 7593 59866
rect 7605 59814 7657 59866
rect 7669 59814 7721 59866
rect 7733 59814 7785 59866
rect 1676 59712 1728 59764
rect 2872 59712 2924 59764
rect 3148 59712 3200 59764
rect 940 59644 992 59696
rect 1492 59576 1544 59628
rect 1400 59508 1452 59560
rect 848 59372 900 59424
rect 2582 59270 2634 59322
rect 2646 59270 2698 59322
rect 2710 59270 2762 59322
rect 2774 59270 2826 59322
rect 2838 59270 2890 59322
rect 5845 59270 5897 59322
rect 5909 59270 5961 59322
rect 5973 59270 6025 59322
rect 6037 59270 6089 59322
rect 6101 59270 6153 59322
rect 9109 59270 9161 59322
rect 9173 59270 9225 59322
rect 9237 59270 9289 59322
rect 9301 59270 9353 59322
rect 9365 59270 9417 59322
rect 9864 59168 9916 59220
rect 756 58964 808 59016
rect 1860 59032 1912 59084
rect 10140 59007 10192 59016
rect 10140 58973 10149 59007
rect 10149 58973 10183 59007
rect 10183 58973 10192 59007
rect 10140 58964 10192 58973
rect 1492 58871 1544 58880
rect 1492 58837 1501 58871
rect 1501 58837 1535 58871
rect 1535 58837 1544 58871
rect 1492 58828 1544 58837
rect 4213 58726 4265 58778
rect 4277 58726 4329 58778
rect 4341 58726 4393 58778
rect 4405 58726 4457 58778
rect 4469 58726 4521 58778
rect 7477 58726 7529 58778
rect 7541 58726 7593 58778
rect 7605 58726 7657 58778
rect 7669 58726 7721 58778
rect 7733 58726 7785 58778
rect 848 58488 900 58540
rect 10140 58531 10192 58540
rect 10140 58497 10149 58531
rect 10149 58497 10183 58531
rect 10183 58497 10192 58531
rect 10140 58488 10192 58497
rect 1400 58284 1452 58336
rect 9956 58327 10008 58336
rect 9956 58293 9965 58327
rect 9965 58293 9999 58327
rect 9999 58293 10008 58327
rect 9956 58284 10008 58293
rect 2582 58182 2634 58234
rect 2646 58182 2698 58234
rect 2710 58182 2762 58234
rect 2774 58182 2826 58234
rect 2838 58182 2890 58234
rect 5845 58182 5897 58234
rect 5909 58182 5961 58234
rect 5973 58182 6025 58234
rect 6037 58182 6089 58234
rect 6101 58182 6153 58234
rect 9109 58182 9161 58234
rect 9173 58182 9225 58234
rect 9237 58182 9289 58234
rect 9301 58182 9353 58234
rect 9365 58182 9417 58234
rect 1860 58012 1912 58064
rect 2872 58012 2924 58064
rect 1492 57944 1544 57996
rect 1952 57876 2004 57928
rect 4712 57876 4764 57928
rect 10140 57919 10192 57928
rect 10140 57885 10149 57919
rect 10149 57885 10183 57919
rect 10183 57885 10192 57919
rect 10140 57876 10192 57885
rect 1124 57740 1176 57792
rect 1308 57740 1360 57792
rect 2136 57740 2188 57792
rect 2780 57740 2832 57792
rect 4213 57638 4265 57690
rect 4277 57638 4329 57690
rect 4341 57638 4393 57690
rect 4405 57638 4457 57690
rect 4469 57638 4521 57690
rect 7477 57638 7529 57690
rect 7541 57638 7593 57690
rect 7605 57638 7657 57690
rect 7669 57638 7721 57690
rect 7733 57638 7785 57690
rect 1676 57536 1728 57588
rect 2136 57536 2188 57588
rect 2412 57536 2464 57588
rect 7196 57536 7248 57588
rect 1124 57468 1176 57520
rect 1492 57400 1544 57452
rect 1952 57400 2004 57452
rect 2320 57400 2372 57452
rect 3332 57400 3384 57452
rect 9956 57332 10008 57384
rect 3700 57264 3752 57316
rect 1676 57196 1728 57248
rect 5448 57196 5500 57248
rect 2582 57094 2634 57146
rect 2646 57094 2698 57146
rect 2710 57094 2762 57146
rect 2774 57094 2826 57146
rect 2838 57094 2890 57146
rect 5845 57094 5897 57146
rect 5909 57094 5961 57146
rect 5973 57094 6025 57146
rect 6037 57094 6089 57146
rect 6101 57094 6153 57146
rect 9109 57094 9161 57146
rect 9173 57094 9225 57146
rect 9237 57094 9289 57146
rect 9301 57094 9353 57146
rect 9365 57094 9417 57146
rect 2320 56924 2372 56976
rect 2596 56856 2648 56908
rect 1676 56831 1728 56840
rect 1676 56797 1685 56831
rect 1685 56797 1719 56831
rect 1719 56797 1728 56831
rect 1676 56788 1728 56797
rect 2780 56924 2832 56976
rect 3332 56924 3384 56976
rect 10140 56831 10192 56840
rect 10140 56797 10149 56831
rect 10149 56797 10183 56831
rect 10183 56797 10192 56831
rect 10140 56788 10192 56797
rect 2504 56763 2556 56772
rect 2504 56729 2513 56763
rect 2513 56729 2547 56763
rect 2547 56729 2556 56763
rect 2504 56720 2556 56729
rect 1492 56695 1544 56704
rect 1492 56661 1501 56695
rect 1501 56661 1535 56695
rect 1535 56661 1544 56695
rect 1492 56652 1544 56661
rect 8760 56652 8812 56704
rect 4213 56550 4265 56602
rect 4277 56550 4329 56602
rect 4341 56550 4393 56602
rect 4405 56550 4457 56602
rect 4469 56550 4521 56602
rect 7477 56550 7529 56602
rect 7541 56550 7593 56602
rect 7605 56550 7657 56602
rect 7669 56550 7721 56602
rect 7733 56550 7785 56602
rect 1400 56448 1452 56500
rect 1676 56448 1728 56500
rect 3608 56448 3660 56500
rect 1860 56380 1912 56432
rect 2320 56380 2372 56432
rect 2780 56380 2832 56432
rect 8852 56312 8904 56364
rect 10140 56355 10192 56364
rect 10140 56321 10149 56355
rect 10149 56321 10183 56355
rect 10183 56321 10192 56355
rect 10140 56312 10192 56321
rect 3240 56244 3292 56296
rect 3608 56244 3660 56296
rect 3976 56244 4028 56296
rect 1860 56176 1912 56228
rect 2872 56176 2924 56228
rect 3056 56176 3108 56228
rect 3148 56151 3200 56160
rect 3148 56117 3157 56151
rect 3157 56117 3191 56151
rect 3191 56117 3200 56151
rect 3148 56108 3200 56117
rect 9956 56151 10008 56160
rect 9956 56117 9965 56151
rect 9965 56117 9999 56151
rect 9999 56117 10008 56151
rect 9956 56108 10008 56117
rect 2582 56006 2634 56058
rect 2646 56006 2698 56058
rect 2710 56006 2762 56058
rect 2774 56006 2826 56058
rect 2838 56006 2890 56058
rect 5845 56006 5897 56058
rect 5909 56006 5961 56058
rect 5973 56006 6025 56058
rect 6037 56006 6089 56058
rect 6101 56006 6153 56058
rect 9109 56006 9161 56058
rect 9173 56006 9225 56058
rect 9237 56006 9289 56058
rect 9301 56006 9353 56058
rect 9365 56006 9417 56058
rect 2412 55904 2464 55956
rect 3332 55836 3384 55888
rect 7932 55768 7984 55820
rect 8668 55700 8720 55752
rect 1492 55607 1544 55616
rect 1492 55573 1501 55607
rect 1501 55573 1535 55607
rect 1535 55573 1544 55607
rect 1492 55564 1544 55573
rect 3148 55632 3200 55684
rect 2504 55564 2556 55616
rect 2780 55564 2832 55616
rect 3976 55607 4028 55616
rect 3976 55573 3985 55607
rect 3985 55573 4019 55607
rect 4019 55573 4028 55607
rect 3976 55564 4028 55573
rect 4213 55462 4265 55514
rect 4277 55462 4329 55514
rect 4341 55462 4393 55514
rect 4405 55462 4457 55514
rect 4469 55462 4521 55514
rect 7477 55462 7529 55514
rect 7541 55462 7593 55514
rect 7605 55462 7657 55514
rect 7669 55462 7721 55514
rect 7733 55462 7785 55514
rect 9956 55360 10008 55412
rect 2780 55292 2832 55344
rect 3240 55292 3292 55344
rect 3976 55292 4028 55344
rect 1860 55267 1912 55276
rect 1860 55233 1863 55267
rect 1863 55233 1912 55267
rect 1860 55224 1912 55233
rect 8392 55224 8444 55276
rect 10140 55267 10192 55276
rect 10140 55233 10149 55267
rect 10149 55233 10183 55267
rect 10183 55233 10192 55267
rect 10140 55224 10192 55233
rect 1676 55156 1728 55208
rect 2780 55088 2832 55140
rect 1676 55020 1728 55072
rect 9956 55063 10008 55072
rect 9956 55029 9965 55063
rect 9965 55029 9999 55063
rect 9999 55029 10008 55063
rect 9956 55020 10008 55029
rect 2582 54918 2634 54970
rect 2646 54918 2698 54970
rect 2710 54918 2762 54970
rect 2774 54918 2826 54970
rect 2838 54918 2890 54970
rect 5845 54918 5897 54970
rect 5909 54918 5961 54970
rect 5973 54918 6025 54970
rect 6037 54918 6089 54970
rect 6101 54918 6153 54970
rect 9109 54918 9161 54970
rect 9173 54918 9225 54970
rect 9237 54918 9289 54970
rect 9301 54918 9353 54970
rect 9365 54918 9417 54970
rect 6828 54612 6880 54664
rect 10140 54655 10192 54664
rect 10140 54621 10149 54655
rect 10149 54621 10183 54655
rect 10183 54621 10192 54655
rect 10140 54612 10192 54621
rect 7288 54544 7340 54596
rect 1492 54519 1544 54528
rect 1492 54485 1501 54519
rect 1501 54485 1535 54519
rect 1535 54485 1544 54519
rect 1492 54476 1544 54485
rect 2228 54519 2280 54528
rect 2228 54485 2237 54519
rect 2237 54485 2271 54519
rect 2271 54485 2280 54519
rect 2228 54476 2280 54485
rect 4213 54374 4265 54426
rect 4277 54374 4329 54426
rect 4341 54374 4393 54426
rect 4405 54374 4457 54426
rect 4469 54374 4521 54426
rect 7477 54374 7529 54426
rect 7541 54374 7593 54426
rect 7605 54374 7657 54426
rect 7669 54374 7721 54426
rect 7733 54374 7785 54426
rect 3056 54272 3108 54324
rect 2504 54136 2556 54188
rect 2964 54136 3016 54188
rect 3332 54136 3384 54188
rect 5724 54136 5776 54188
rect 6276 54136 6328 54188
rect 9772 54136 9824 54188
rect 1676 54068 1728 54120
rect 10048 53975 10100 53984
rect 10048 53941 10057 53975
rect 10057 53941 10091 53975
rect 10091 53941 10100 53975
rect 10048 53932 10100 53941
rect 2582 53830 2634 53882
rect 2646 53830 2698 53882
rect 2710 53830 2762 53882
rect 2774 53830 2826 53882
rect 2838 53830 2890 53882
rect 5845 53830 5897 53882
rect 5909 53830 5961 53882
rect 5973 53830 6025 53882
rect 6037 53830 6089 53882
rect 6101 53830 6153 53882
rect 9109 53830 9161 53882
rect 9173 53830 9225 53882
rect 9237 53830 9289 53882
rect 9301 53830 9353 53882
rect 9365 53830 9417 53882
rect 1768 53660 1820 53712
rect 1492 53524 1544 53576
rect 1860 53567 1912 53576
rect 1860 53533 1863 53567
rect 1863 53533 1912 53567
rect 1860 53524 1912 53533
rect 8024 53524 8076 53576
rect 9956 53456 10008 53508
rect 1768 53388 1820 53440
rect 2136 53388 2188 53440
rect 2780 53388 2832 53440
rect 4213 53286 4265 53338
rect 4277 53286 4329 53338
rect 4341 53286 4393 53338
rect 4405 53286 4457 53338
rect 4469 53286 4521 53338
rect 7477 53286 7529 53338
rect 7541 53286 7593 53338
rect 7605 53286 7657 53338
rect 7669 53286 7721 53338
rect 7733 53286 7785 53338
rect 1492 53184 1544 53236
rect 1676 53184 1728 53236
rect 2504 53184 2556 53236
rect 6644 53116 6696 53168
rect 8116 53048 8168 53100
rect 9864 53091 9916 53100
rect 9864 53057 9873 53091
rect 9873 53057 9907 53091
rect 9907 53057 9916 53091
rect 9864 53048 9916 53057
rect 5264 52980 5316 53032
rect 3056 52955 3108 52964
rect 3056 52921 3065 52955
rect 3065 52921 3099 52955
rect 3099 52921 3108 52955
rect 3056 52912 3108 52921
rect 1400 52844 1452 52896
rect 2228 52887 2280 52896
rect 2228 52853 2237 52887
rect 2237 52853 2271 52887
rect 2271 52853 2280 52887
rect 2228 52844 2280 52853
rect 10048 52887 10100 52896
rect 10048 52853 10057 52887
rect 10057 52853 10091 52887
rect 10091 52853 10100 52887
rect 10048 52844 10100 52853
rect 2582 52742 2634 52794
rect 2646 52742 2698 52794
rect 2710 52742 2762 52794
rect 2774 52742 2826 52794
rect 2838 52742 2890 52794
rect 5845 52742 5897 52794
rect 5909 52742 5961 52794
rect 5973 52742 6025 52794
rect 6037 52742 6089 52794
rect 6101 52742 6153 52794
rect 9109 52742 9161 52794
rect 9173 52742 9225 52794
rect 9237 52742 9289 52794
rect 9301 52742 9353 52794
rect 9365 52742 9417 52794
rect 2412 52640 2464 52692
rect 9772 52640 9824 52692
rect 1216 52436 1268 52488
rect 2228 52436 2280 52488
rect 2412 52436 2464 52488
rect 3056 52436 3108 52488
rect 2872 52368 2924 52420
rect 3148 52368 3200 52420
rect 1492 52343 1544 52352
rect 1492 52309 1501 52343
rect 1501 52309 1535 52343
rect 1535 52309 1544 52343
rect 1492 52300 1544 52309
rect 2320 52300 2372 52352
rect 7380 52300 7432 52352
rect 10048 52343 10100 52352
rect 10048 52309 10057 52343
rect 10057 52309 10091 52343
rect 10091 52309 10100 52343
rect 10048 52300 10100 52309
rect 4213 52198 4265 52250
rect 4277 52198 4329 52250
rect 4341 52198 4393 52250
rect 4405 52198 4457 52250
rect 4469 52198 4521 52250
rect 7477 52198 7529 52250
rect 7541 52198 7593 52250
rect 7605 52198 7657 52250
rect 7669 52198 7721 52250
rect 7733 52198 7785 52250
rect 3148 52096 3200 52148
rect 9864 52096 9916 52148
rect 572 52028 624 52080
rect 2320 51960 2372 52012
rect 2964 51960 3016 52012
rect 3056 52003 3108 52012
rect 3056 51969 3077 52003
rect 3077 51969 3108 52003
rect 3056 51960 3108 51969
rect 2136 51824 2188 51876
rect 2320 51824 2372 51876
rect 2872 51824 2924 51876
rect 3148 51824 3200 51876
rect 1308 51756 1360 51808
rect 1676 51756 1728 51808
rect 8208 51756 8260 51808
rect 2582 51654 2634 51706
rect 2646 51654 2698 51706
rect 2710 51654 2762 51706
rect 2774 51654 2826 51706
rect 2838 51654 2890 51706
rect 5845 51654 5897 51706
rect 5909 51654 5961 51706
rect 5973 51654 6025 51706
rect 6037 51654 6089 51706
rect 6101 51654 6153 51706
rect 9109 51654 9161 51706
rect 9173 51654 9225 51706
rect 9237 51654 9289 51706
rect 9301 51654 9353 51706
rect 9365 51654 9417 51706
rect 3792 51552 3844 51604
rect 1676 51391 1728 51400
rect 1676 51357 1685 51391
rect 1685 51357 1719 51391
rect 1719 51357 1728 51391
rect 1676 51348 1728 51357
rect 2412 51484 2464 51536
rect 2688 51484 2740 51536
rect 3700 51484 3752 51536
rect 2780 51348 2832 51400
rect 3148 51416 3200 51468
rect 3056 51391 3108 51400
rect 3056 51357 3065 51391
rect 3065 51357 3099 51391
rect 3099 51357 3108 51391
rect 3056 51348 3108 51357
rect 9864 51391 9916 51400
rect 9864 51357 9873 51391
rect 9873 51357 9907 51391
rect 9907 51357 9916 51391
rect 9864 51348 9916 51357
rect 2964 51280 3016 51332
rect 1400 51212 1452 51264
rect 1676 51212 1728 51264
rect 2228 51255 2280 51264
rect 2228 51221 2237 51255
rect 2237 51221 2271 51255
rect 2271 51221 2280 51255
rect 2228 51212 2280 51221
rect 10048 51255 10100 51264
rect 10048 51221 10057 51255
rect 10057 51221 10091 51255
rect 10091 51221 10100 51255
rect 10048 51212 10100 51221
rect 4213 51110 4265 51162
rect 4277 51110 4329 51162
rect 4341 51110 4393 51162
rect 4405 51110 4457 51162
rect 4469 51110 4521 51162
rect 7477 51110 7529 51162
rect 7541 51110 7593 51162
rect 7605 51110 7657 51162
rect 7669 51110 7721 51162
rect 7733 51110 7785 51162
rect 2228 51051 2280 51060
rect 2228 51017 2237 51051
rect 2237 51017 2271 51051
rect 2271 51017 2280 51051
rect 2228 51008 2280 51017
rect 3240 51008 3292 51060
rect 2228 50872 2280 50924
rect 2504 50872 2556 50924
rect 3056 50940 3108 50992
rect 3700 51008 3752 51060
rect 2780 50915 2832 50924
rect 2780 50881 2789 50915
rect 2789 50881 2823 50915
rect 2823 50881 2832 50915
rect 2780 50872 2832 50881
rect 3056 50804 3108 50856
rect 204 50736 256 50788
rect 1492 50711 1544 50720
rect 1492 50677 1501 50711
rect 1501 50677 1535 50711
rect 1535 50677 1544 50711
rect 1492 50668 1544 50677
rect 1952 50736 2004 50788
rect 2688 50736 2740 50788
rect 3700 50872 3752 50924
rect 10048 50711 10100 50720
rect 10048 50677 10057 50711
rect 10057 50677 10091 50711
rect 10091 50677 10100 50711
rect 10048 50668 10100 50677
rect 2582 50566 2634 50618
rect 2646 50566 2698 50618
rect 2710 50566 2762 50618
rect 2774 50566 2826 50618
rect 2838 50566 2890 50618
rect 5845 50566 5897 50618
rect 5909 50566 5961 50618
rect 5973 50566 6025 50618
rect 6037 50566 6089 50618
rect 6101 50566 6153 50618
rect 9109 50566 9161 50618
rect 9173 50566 9225 50618
rect 9237 50566 9289 50618
rect 9301 50566 9353 50618
rect 9365 50566 9417 50618
rect 112 50464 164 50516
rect 1676 50464 1728 50516
rect 3240 50464 3292 50516
rect 2412 50396 2464 50448
rect 9864 50464 9916 50516
rect 1676 50328 1728 50380
rect 3056 50328 3108 50380
rect 1584 50303 1636 50312
rect 1584 50269 1593 50303
rect 1593 50269 1627 50303
rect 1627 50269 1636 50303
rect 1584 50260 1636 50269
rect 1860 50260 1912 50312
rect 2228 50260 2280 50312
rect 3240 50260 3292 50312
rect 3884 50260 3936 50312
rect 1216 50192 1268 50244
rect 2780 50192 2832 50244
rect 3056 50192 3108 50244
rect 3424 50192 3476 50244
rect 1584 50124 1636 50176
rect 3240 50124 3292 50176
rect 3700 50124 3752 50176
rect 10968 50371 11020 50380
rect 10968 50337 10977 50371
rect 10977 50337 11011 50371
rect 11011 50337 11020 50371
rect 10968 50328 11020 50337
rect 10048 50167 10100 50176
rect 10048 50133 10057 50167
rect 10057 50133 10091 50167
rect 10091 50133 10100 50167
rect 10048 50124 10100 50133
rect 4213 50022 4265 50074
rect 4277 50022 4329 50074
rect 4341 50022 4393 50074
rect 4405 50022 4457 50074
rect 4469 50022 4521 50074
rect 7477 50022 7529 50074
rect 7541 50022 7593 50074
rect 7605 50022 7657 50074
rect 7669 50022 7721 50074
rect 7733 50022 7785 50074
rect 1768 49920 1820 49972
rect 2780 49920 2832 49972
rect 2228 49784 2280 49836
rect 2412 49827 2464 49836
rect 2412 49793 2421 49827
rect 2421 49793 2455 49827
rect 2455 49793 2464 49827
rect 2412 49784 2464 49793
rect 296 49716 348 49768
rect 1676 49716 1728 49768
rect 2412 49580 2464 49632
rect 4160 49852 4212 49904
rect 4896 49852 4948 49904
rect 3700 49784 3752 49836
rect 3884 49784 3936 49836
rect 10968 49784 11020 49836
rect 9680 49716 9732 49768
rect 2582 49478 2634 49530
rect 2646 49478 2698 49530
rect 2710 49478 2762 49530
rect 2774 49478 2826 49530
rect 2838 49478 2890 49530
rect 5845 49478 5897 49530
rect 5909 49478 5961 49530
rect 5973 49478 6025 49530
rect 6037 49478 6089 49530
rect 6101 49478 6153 49530
rect 9109 49478 9161 49530
rect 9173 49478 9225 49530
rect 9237 49478 9289 49530
rect 9301 49478 9353 49530
rect 9365 49478 9417 49530
rect 664 49376 716 49428
rect 1584 49376 1636 49428
rect 1768 49376 1820 49428
rect 1952 49376 2004 49428
rect 4804 49376 4856 49428
rect 5172 49376 5224 49428
rect 1400 49172 1452 49224
rect 2228 49308 2280 49360
rect 1952 49215 2004 49224
rect 1952 49181 1961 49215
rect 1961 49181 1995 49215
rect 1995 49181 2004 49215
rect 1952 49172 2004 49181
rect 2688 49215 2740 49224
rect 2688 49181 2697 49215
rect 2697 49181 2731 49215
rect 2731 49181 2740 49215
rect 2688 49172 2740 49181
rect 3884 49240 3936 49292
rect 5172 49240 5224 49292
rect 3700 49104 3752 49156
rect 9588 49172 9640 49224
rect 1400 49079 1452 49088
rect 1400 49045 1409 49079
rect 1409 49045 1443 49079
rect 1443 49045 1452 49079
rect 1400 49036 1452 49045
rect 2780 49036 2832 49088
rect 9864 49036 9916 49088
rect 10048 49079 10100 49088
rect 10048 49045 10057 49079
rect 10057 49045 10091 49079
rect 10091 49045 10100 49079
rect 10048 49036 10100 49045
rect 4213 48934 4265 48986
rect 4277 48934 4329 48986
rect 4341 48934 4393 48986
rect 4405 48934 4457 48986
rect 4469 48934 4521 48986
rect 7477 48934 7529 48986
rect 7541 48934 7593 48986
rect 7605 48934 7657 48986
rect 7669 48934 7721 48986
rect 7733 48934 7785 48986
rect 2228 48875 2280 48884
rect 2228 48841 2237 48875
rect 2237 48841 2271 48875
rect 2271 48841 2280 48875
rect 2228 48832 2280 48841
rect 2688 48832 2740 48884
rect 6460 48832 6512 48884
rect 664 48764 716 48816
rect 1952 48764 2004 48816
rect 2228 48696 2280 48748
rect 1492 48535 1544 48544
rect 1492 48501 1501 48535
rect 1501 48501 1535 48535
rect 1535 48501 1544 48535
rect 1492 48492 1544 48501
rect 3700 48696 3752 48748
rect 9772 48696 9824 48748
rect 6092 48560 6144 48612
rect 5724 48492 5776 48544
rect 6184 48492 6236 48544
rect 10048 48535 10100 48544
rect 10048 48501 10057 48535
rect 10057 48501 10091 48535
rect 10091 48501 10100 48535
rect 10048 48492 10100 48501
rect 2582 48390 2634 48442
rect 2646 48390 2698 48442
rect 2710 48390 2762 48442
rect 2774 48390 2826 48442
rect 2838 48390 2890 48442
rect 5845 48390 5897 48442
rect 5909 48390 5961 48442
rect 5973 48390 6025 48442
rect 6037 48390 6089 48442
rect 6101 48390 6153 48442
rect 9109 48390 9161 48442
rect 9173 48390 9225 48442
rect 9237 48390 9289 48442
rect 9301 48390 9353 48442
rect 9365 48390 9417 48442
rect 388 48288 440 48340
rect 2412 48288 2464 48340
rect 4620 48288 4672 48340
rect 2688 48220 2740 48272
rect 204 48152 256 48204
rect 2044 48084 2096 48136
rect 5080 48152 5132 48204
rect 9772 48220 9824 48272
rect 388 48016 440 48068
rect 1492 47991 1544 48000
rect 1492 47957 1501 47991
rect 1501 47957 1535 47991
rect 1535 47957 1544 47991
rect 1492 47948 1544 47957
rect 1768 48016 1820 48068
rect 3240 48084 3292 48136
rect 3148 47948 3200 48000
rect 4213 47846 4265 47898
rect 4277 47846 4329 47898
rect 4341 47846 4393 47898
rect 4405 47846 4457 47898
rect 4469 47846 4521 47898
rect 7477 47846 7529 47898
rect 7541 47846 7593 47898
rect 7605 47846 7657 47898
rect 7669 47846 7721 47898
rect 7733 47846 7785 47898
rect 2964 47744 3016 47796
rect 2044 47676 2096 47728
rect 6184 47676 6236 47728
rect 3148 47608 3200 47660
rect 9680 47608 9732 47660
rect 7932 47540 7984 47592
rect 9036 47472 9088 47524
rect 10048 47515 10100 47524
rect 10048 47481 10057 47515
rect 10057 47481 10091 47515
rect 10091 47481 10100 47515
rect 10048 47472 10100 47481
rect 1492 47447 1544 47456
rect 1492 47413 1501 47447
rect 1501 47413 1535 47447
rect 1535 47413 1544 47447
rect 1492 47404 1544 47413
rect 2228 47447 2280 47456
rect 2228 47413 2237 47447
rect 2237 47413 2271 47447
rect 2271 47413 2280 47447
rect 2228 47404 2280 47413
rect 2582 47302 2634 47354
rect 2646 47302 2698 47354
rect 2710 47302 2762 47354
rect 2774 47302 2826 47354
rect 2838 47302 2890 47354
rect 5845 47302 5897 47354
rect 5909 47302 5961 47354
rect 5973 47302 6025 47354
rect 6037 47302 6089 47354
rect 6101 47302 6153 47354
rect 9109 47302 9161 47354
rect 9173 47302 9225 47354
rect 9237 47302 9289 47354
rect 9301 47302 9353 47354
rect 9365 47302 9417 47354
rect 2320 47200 2372 47252
rect 3792 47200 3844 47252
rect 4620 47132 4672 47184
rect 4804 47132 4856 47184
rect 8944 47064 8996 47116
rect 2320 47039 2372 47048
rect 2320 47005 2329 47039
rect 2329 47005 2363 47039
rect 2363 47005 2372 47039
rect 2320 46996 2372 47005
rect 4804 46996 4856 47048
rect 1492 46903 1544 46912
rect 1492 46869 1501 46903
rect 1501 46869 1535 46903
rect 1535 46869 1544 46903
rect 1492 46860 1544 46869
rect 2964 46860 3016 46912
rect 10048 46903 10100 46912
rect 10048 46869 10057 46903
rect 10057 46869 10091 46903
rect 10091 46869 10100 46903
rect 10048 46860 10100 46869
rect 4213 46758 4265 46810
rect 4277 46758 4329 46810
rect 4341 46758 4393 46810
rect 4405 46758 4457 46810
rect 4469 46758 4521 46810
rect 7477 46758 7529 46810
rect 7541 46758 7593 46810
rect 7605 46758 7657 46810
rect 7669 46758 7721 46810
rect 7733 46758 7785 46810
rect 1952 46656 2004 46708
rect 2412 46656 2464 46708
rect 2596 46656 2648 46708
rect 9588 46656 9640 46708
rect 1492 46359 1544 46368
rect 1492 46325 1501 46359
rect 1501 46325 1535 46359
rect 1535 46325 1544 46359
rect 1492 46316 1544 46325
rect 2596 46520 2648 46572
rect 2964 46520 3016 46572
rect 3240 46520 3292 46572
rect 3884 46520 3936 46572
rect 9864 46563 9916 46572
rect 9864 46529 9873 46563
rect 9873 46529 9907 46563
rect 9907 46529 9916 46563
rect 9864 46520 9916 46529
rect 3240 46384 3292 46436
rect 4712 46384 4764 46436
rect 5172 46384 5224 46436
rect 4620 46316 4672 46368
rect 10048 46359 10100 46368
rect 10048 46325 10057 46359
rect 10057 46325 10091 46359
rect 10091 46325 10100 46359
rect 10048 46316 10100 46325
rect 2582 46214 2634 46266
rect 2646 46214 2698 46266
rect 2710 46214 2762 46266
rect 2774 46214 2826 46266
rect 2838 46214 2890 46266
rect 5845 46214 5897 46266
rect 5909 46214 5961 46266
rect 5973 46214 6025 46266
rect 6037 46214 6089 46266
rect 6101 46214 6153 46266
rect 9109 46214 9161 46266
rect 9173 46214 9225 46266
rect 9237 46214 9289 46266
rect 9301 46214 9353 46266
rect 9365 46214 9417 46266
rect 1860 46112 1912 46164
rect 2136 46112 2188 46164
rect 4712 46044 4764 46096
rect 5264 46044 5316 46096
rect 5724 46044 5776 46096
rect 6644 46044 6696 46096
rect 480 45976 532 46028
rect 4896 45976 4948 46028
rect 5448 45976 5500 46028
rect 1768 45951 1820 45960
rect 1768 45917 1777 45951
rect 1777 45917 1811 45951
rect 1811 45917 1820 45951
rect 1768 45908 1820 45917
rect 2136 45908 2188 45960
rect 2320 45908 2372 45960
rect 4528 45840 4580 45892
rect 5448 45840 5500 45892
rect 7840 46112 7892 46164
rect 7288 46044 7340 46096
rect 7380 46044 7432 46096
rect 7932 46044 7984 46096
rect 1952 45772 2004 45824
rect 2412 45772 2464 45824
rect 2964 45772 3016 45824
rect 7104 45772 7156 45824
rect 7196 45772 7248 45824
rect 4213 45670 4265 45722
rect 4277 45670 4329 45722
rect 4341 45670 4393 45722
rect 4405 45670 4457 45722
rect 4469 45670 4521 45722
rect 7477 45670 7529 45722
rect 7541 45670 7593 45722
rect 7605 45670 7657 45722
rect 7669 45670 7721 45722
rect 7733 45670 7785 45722
rect 7932 45432 7984 45484
rect 3424 45407 3476 45416
rect 3424 45373 3433 45407
rect 3433 45373 3467 45407
rect 3467 45373 3476 45407
rect 3424 45364 3476 45373
rect 3700 45407 3752 45416
rect 3700 45373 3709 45407
rect 3709 45373 3743 45407
rect 3743 45373 3752 45407
rect 3700 45364 3752 45373
rect 1492 45271 1544 45280
rect 1492 45237 1501 45271
rect 1501 45237 1535 45271
rect 1535 45237 1544 45271
rect 1492 45228 1544 45237
rect 10048 45271 10100 45280
rect 10048 45237 10057 45271
rect 10057 45237 10091 45271
rect 10091 45237 10100 45271
rect 10048 45228 10100 45237
rect 2582 45126 2634 45178
rect 2646 45126 2698 45178
rect 2710 45126 2762 45178
rect 2774 45126 2826 45178
rect 2838 45126 2890 45178
rect 5845 45126 5897 45178
rect 5909 45126 5961 45178
rect 5973 45126 6025 45178
rect 6037 45126 6089 45178
rect 6101 45126 6153 45178
rect 9109 45126 9161 45178
rect 9173 45126 9225 45178
rect 9237 45126 9289 45178
rect 9301 45126 9353 45178
rect 9365 45126 9417 45178
rect 1032 44888 1084 44940
rect 1768 44820 1820 44872
rect 2044 44888 2096 44940
rect 2412 44888 2464 44940
rect 2964 44820 3016 44872
rect 2412 44727 2464 44736
rect 2412 44693 2421 44727
rect 2421 44693 2455 44727
rect 2455 44693 2464 44727
rect 2412 44684 2464 44693
rect 3700 44820 3752 44872
rect 3792 44863 3844 44872
rect 3792 44829 3801 44863
rect 3801 44829 3835 44863
rect 3835 44829 3844 44863
rect 3792 44820 3844 44829
rect 5080 44820 5132 44872
rect 3240 44684 3292 44736
rect 3700 44684 3752 44736
rect 9864 44684 9916 44736
rect 10048 44727 10100 44736
rect 10048 44693 10057 44727
rect 10057 44693 10091 44727
rect 10091 44693 10100 44727
rect 10048 44684 10100 44693
rect 4213 44582 4265 44634
rect 4277 44582 4329 44634
rect 4341 44582 4393 44634
rect 4405 44582 4457 44634
rect 4469 44582 4521 44634
rect 7477 44582 7529 44634
rect 7541 44582 7593 44634
rect 7605 44582 7657 44634
rect 7669 44582 7721 44634
rect 7733 44582 7785 44634
rect 1124 44480 1176 44532
rect 1768 44344 1820 44396
rect 3332 44480 3384 44532
rect 3608 44480 3660 44532
rect 3056 44387 3108 44396
rect 3056 44353 3065 44387
rect 3065 44353 3099 44387
rect 3099 44353 3108 44387
rect 3056 44344 3108 44353
rect 3240 44387 3292 44396
rect 3240 44353 3249 44387
rect 3249 44353 3283 44387
rect 3283 44353 3292 44387
rect 3240 44344 3292 44353
rect 3332 44276 3384 44328
rect 3792 44344 3844 44396
rect 4436 44344 4488 44396
rect 5264 44276 5316 44328
rect 664 44140 716 44192
rect 1124 44140 1176 44192
rect 2412 44140 2464 44192
rect 3884 44208 3936 44260
rect 4436 44208 4488 44260
rect 5448 44140 5500 44192
rect 112 44004 164 44056
rect 664 44004 716 44056
rect 2582 44038 2634 44090
rect 2646 44038 2698 44090
rect 2710 44038 2762 44090
rect 2774 44038 2826 44090
rect 2838 44038 2890 44090
rect 5845 44038 5897 44090
rect 5909 44038 5961 44090
rect 5973 44038 6025 44090
rect 6037 44038 6089 44090
rect 6101 44038 6153 44090
rect 9109 44038 9161 44090
rect 9173 44038 9225 44090
rect 9237 44038 9289 44090
rect 9301 44038 9353 44090
rect 9365 44038 9417 44090
rect 1584 43979 1636 43988
rect 1584 43945 1593 43979
rect 1593 43945 1627 43979
rect 1627 43945 1636 43979
rect 1584 43936 1636 43945
rect 1400 43775 1452 43784
rect 1400 43741 1409 43775
rect 1409 43741 1443 43775
rect 1443 43741 1452 43775
rect 1400 43732 1452 43741
rect 2228 43732 2280 43784
rect 8300 43936 8352 43988
rect 4436 43911 4488 43920
rect 4436 43877 4445 43911
rect 4445 43877 4479 43911
rect 4479 43877 4488 43911
rect 4436 43868 4488 43877
rect 3608 43800 3660 43852
rect 3424 43732 3476 43784
rect 5080 43775 5132 43784
rect 1768 43664 1820 43716
rect 5080 43741 5089 43775
rect 5089 43741 5123 43775
rect 5123 43741 5132 43775
rect 5080 43732 5132 43741
rect 9864 43775 9916 43784
rect 9864 43741 9873 43775
rect 9873 43741 9907 43775
rect 9907 43741 9916 43775
rect 9864 43732 9916 43741
rect 5448 43664 5500 43716
rect 2228 43639 2280 43648
rect 2228 43605 2237 43639
rect 2237 43605 2271 43639
rect 2271 43605 2280 43639
rect 2228 43596 2280 43605
rect 3056 43639 3108 43648
rect 3056 43605 3065 43639
rect 3065 43605 3099 43639
rect 3099 43605 3108 43639
rect 3056 43596 3108 43605
rect 9864 43596 9916 43648
rect 10048 43639 10100 43648
rect 10048 43605 10057 43639
rect 10057 43605 10091 43639
rect 10091 43605 10100 43639
rect 10048 43596 10100 43605
rect 4213 43494 4265 43546
rect 4277 43494 4329 43546
rect 4341 43494 4393 43546
rect 4405 43494 4457 43546
rect 4469 43494 4521 43546
rect 7477 43494 7529 43546
rect 7541 43494 7593 43546
rect 7605 43494 7657 43546
rect 7669 43494 7721 43546
rect 7733 43494 7785 43546
rect 940 43392 992 43444
rect 1768 43256 1820 43308
rect 1492 43188 1544 43240
rect 1768 43120 1820 43172
rect 1492 43095 1544 43104
rect 1492 43061 1501 43095
rect 1501 43061 1535 43095
rect 1535 43061 1544 43095
rect 1492 43052 1544 43061
rect 3332 43256 3384 43308
rect 9864 43299 9916 43308
rect 9864 43265 9873 43299
rect 9873 43265 9907 43299
rect 9907 43265 9916 43299
rect 9864 43256 9916 43265
rect 2872 43188 2924 43240
rect 5448 43052 5500 43104
rect 10048 43095 10100 43104
rect 10048 43061 10057 43095
rect 10057 43061 10091 43095
rect 10091 43061 10100 43095
rect 10048 43052 10100 43061
rect 2582 42950 2634 43002
rect 2646 42950 2698 43002
rect 2710 42950 2762 43002
rect 2774 42950 2826 43002
rect 2838 42950 2890 43002
rect 5845 42950 5897 43002
rect 5909 42950 5961 43002
rect 5973 42950 6025 43002
rect 6037 42950 6089 43002
rect 6101 42950 6153 43002
rect 9109 42950 9161 43002
rect 9173 42950 9225 43002
rect 9237 42950 9289 43002
rect 9301 42950 9353 43002
rect 9365 42950 9417 43002
rect 2136 42848 2188 42900
rect 3332 42848 3384 42900
rect 4528 42780 4580 42832
rect 2320 42644 2372 42696
rect 9864 42687 9916 42696
rect 9864 42653 9873 42687
rect 9873 42653 9907 42687
rect 9907 42653 9916 42687
rect 9864 42644 9916 42653
rect 1400 42508 1452 42560
rect 2228 42551 2280 42560
rect 2228 42517 2237 42551
rect 2237 42517 2271 42551
rect 2271 42517 2280 42551
rect 2228 42508 2280 42517
rect 10048 42551 10100 42560
rect 10048 42517 10057 42551
rect 10057 42517 10091 42551
rect 10091 42517 10100 42551
rect 10048 42508 10100 42517
rect 4213 42406 4265 42458
rect 4277 42406 4329 42458
rect 4341 42406 4393 42458
rect 4405 42406 4457 42458
rect 4469 42406 4521 42458
rect 7477 42406 7529 42458
rect 7541 42406 7593 42458
rect 7605 42406 7657 42458
rect 7669 42406 7721 42458
rect 7733 42406 7785 42458
rect 5724 42304 5776 42356
rect 3424 42279 3476 42288
rect 3424 42245 3433 42279
rect 3433 42245 3467 42279
rect 3467 42245 3476 42279
rect 3424 42236 3476 42245
rect 3608 42236 3660 42288
rect 4344 42279 4396 42288
rect 4344 42245 4353 42279
rect 4353 42245 4387 42279
rect 4387 42245 4396 42279
rect 4344 42236 4396 42245
rect 5080 42236 5132 42288
rect 4528 42168 4580 42220
rect 4988 42168 5040 42220
rect 3976 42032 4028 42084
rect 1492 42007 1544 42016
rect 1492 41973 1501 42007
rect 1501 41973 1535 42007
rect 1535 41973 1544 42007
rect 1492 41964 1544 41973
rect 2582 41862 2634 41914
rect 2646 41862 2698 41914
rect 2710 41862 2762 41914
rect 2774 41862 2826 41914
rect 2838 41862 2890 41914
rect 5845 41862 5897 41914
rect 5909 41862 5961 41914
rect 5973 41862 6025 41914
rect 6037 41862 6089 41914
rect 6101 41862 6153 41914
rect 9109 41862 9161 41914
rect 9173 41862 9225 41914
rect 9237 41862 9289 41914
rect 9301 41862 9353 41914
rect 9365 41862 9417 41914
rect 1308 41760 1360 41812
rect 9864 41760 9916 41812
rect 4160 41624 4212 41676
rect 4620 41624 4672 41676
rect 1768 41556 1820 41608
rect 1032 41488 1084 41540
rect 3240 41556 3292 41608
rect 4344 41556 4396 41608
rect 4804 41556 4856 41608
rect 5632 41556 5684 41608
rect 6368 41556 6420 41608
rect 6460 41488 6512 41540
rect 1400 41420 1452 41472
rect 3700 41420 3752 41472
rect 5356 41420 5408 41472
rect 5724 41420 5776 41472
rect 6092 41420 6144 41472
rect 6368 41420 6420 41472
rect 10048 41463 10100 41472
rect 10048 41429 10057 41463
rect 10057 41429 10091 41463
rect 10091 41429 10100 41463
rect 10048 41420 10100 41429
rect 4213 41318 4265 41370
rect 4277 41318 4329 41370
rect 4341 41318 4393 41370
rect 4405 41318 4457 41370
rect 4469 41318 4521 41370
rect 7477 41318 7529 41370
rect 7541 41318 7593 41370
rect 7605 41318 7657 41370
rect 7669 41318 7721 41370
rect 7733 41318 7785 41370
rect 1584 41216 1636 41268
rect 1676 41216 1728 41268
rect 6276 41216 6328 41268
rect 2228 41148 2280 41200
rect 1492 41123 1544 41132
rect 1492 41089 1501 41123
rect 1501 41089 1535 41123
rect 1535 41089 1544 41123
rect 1492 41080 1544 41089
rect 1768 41123 1820 41132
rect 1768 41089 1777 41123
rect 1777 41089 1811 41123
rect 1811 41089 1820 41123
rect 1768 41080 1820 41089
rect 5540 41080 5592 41132
rect 6276 41080 6328 41132
rect 9864 41123 9916 41132
rect 9864 41089 9873 41123
rect 9873 41089 9907 41123
rect 9907 41089 9916 41123
rect 9864 41080 9916 41089
rect 2320 40944 2372 40996
rect 5540 40944 5592 40996
rect 5908 40944 5960 40996
rect 10048 40919 10100 40928
rect 10048 40885 10057 40919
rect 10057 40885 10091 40919
rect 10091 40885 10100 40919
rect 10048 40876 10100 40885
rect 2582 40774 2634 40826
rect 2646 40774 2698 40826
rect 2710 40774 2762 40826
rect 2774 40774 2826 40826
rect 2838 40774 2890 40826
rect 5845 40774 5897 40826
rect 5909 40774 5961 40826
rect 5973 40774 6025 40826
rect 6037 40774 6089 40826
rect 6101 40774 6153 40826
rect 9109 40774 9161 40826
rect 9173 40774 9225 40826
rect 9237 40774 9289 40826
rect 9301 40774 9353 40826
rect 9365 40774 9417 40826
rect 3792 40715 3844 40724
rect 3792 40681 3801 40715
rect 3801 40681 3835 40715
rect 3835 40681 3844 40715
rect 3792 40672 3844 40681
rect 3332 40604 3384 40656
rect 3516 40604 3568 40656
rect 2780 40536 2832 40588
rect 3056 40536 3108 40588
rect 1676 40511 1728 40520
rect 1676 40477 1685 40511
rect 1685 40477 1719 40511
rect 1719 40477 1728 40511
rect 1676 40468 1728 40477
rect 3516 40468 3568 40520
rect 1492 40375 1544 40384
rect 1492 40341 1501 40375
rect 1501 40341 1535 40375
rect 1535 40341 1544 40375
rect 1492 40332 1544 40341
rect 1676 40332 1728 40384
rect 1860 40332 1912 40384
rect 2320 40375 2372 40384
rect 2320 40341 2329 40375
rect 2329 40341 2363 40375
rect 2363 40341 2372 40375
rect 2320 40332 2372 40341
rect 3056 40375 3108 40384
rect 3056 40341 3065 40375
rect 3065 40341 3099 40375
rect 3099 40341 3108 40375
rect 3056 40332 3108 40341
rect 3700 40400 3752 40452
rect 4213 40230 4265 40282
rect 4277 40230 4329 40282
rect 4341 40230 4393 40282
rect 4405 40230 4457 40282
rect 4469 40230 4521 40282
rect 7477 40230 7529 40282
rect 7541 40230 7593 40282
rect 7605 40230 7657 40282
rect 7669 40230 7721 40282
rect 7733 40230 7785 40282
rect 756 40128 808 40180
rect 2780 40103 2832 40112
rect 2780 40069 2789 40103
rect 2789 40069 2823 40103
rect 2823 40069 2832 40103
rect 2780 40060 2832 40069
rect 3240 40060 3292 40112
rect 3976 40060 4028 40112
rect 1860 39992 1912 40044
rect 2872 39992 2924 40044
rect 3516 39992 3568 40044
rect 3792 39992 3844 40044
rect 4528 39992 4580 40044
rect 2872 39856 2924 39908
rect 5172 39856 5224 39908
rect 10048 39899 10100 39908
rect 10048 39865 10057 39899
rect 10057 39865 10091 39899
rect 10091 39865 10100 39899
rect 10048 39856 10100 39865
rect 3884 39788 3936 39840
rect 4344 39788 4396 39840
rect 8484 39788 8536 39840
rect 2582 39686 2634 39738
rect 2646 39686 2698 39738
rect 2710 39686 2762 39738
rect 2774 39686 2826 39738
rect 2838 39686 2890 39738
rect 5845 39686 5897 39738
rect 5909 39686 5961 39738
rect 5973 39686 6025 39738
rect 6037 39686 6089 39738
rect 6101 39686 6153 39738
rect 9109 39686 9161 39738
rect 9173 39686 9225 39738
rect 9237 39686 9289 39738
rect 9301 39686 9353 39738
rect 9365 39686 9417 39738
rect 4896 39584 4948 39636
rect 5172 39516 5224 39568
rect 2412 39423 2464 39432
rect 2412 39389 2421 39423
rect 2421 39389 2455 39423
rect 2455 39389 2464 39423
rect 2412 39380 2464 39389
rect 4344 39448 4396 39500
rect 1860 39312 1912 39364
rect 3884 39380 3936 39432
rect 4068 39380 4120 39432
rect 4528 39312 4580 39364
rect 1400 39244 1452 39296
rect 2228 39287 2280 39296
rect 2228 39253 2237 39287
rect 2237 39253 2271 39287
rect 2271 39253 2280 39287
rect 2228 39244 2280 39253
rect 2964 39287 3016 39296
rect 2964 39253 2973 39287
rect 2973 39253 3007 39287
rect 3007 39253 3016 39287
rect 2964 39244 3016 39253
rect 3792 39244 3844 39296
rect 5172 39244 5224 39296
rect 10048 39287 10100 39296
rect 10048 39253 10057 39287
rect 10057 39253 10091 39287
rect 10091 39253 10100 39287
rect 10048 39244 10100 39253
rect 4213 39142 4265 39194
rect 4277 39142 4329 39194
rect 4341 39142 4393 39194
rect 4405 39142 4457 39194
rect 4469 39142 4521 39194
rect 7477 39142 7529 39194
rect 7541 39142 7593 39194
rect 7605 39142 7657 39194
rect 7669 39142 7721 39194
rect 7733 39142 7785 39194
rect 848 38972 900 39024
rect 2412 38972 2464 39024
rect 1860 38947 1912 38956
rect 1860 38913 1869 38947
rect 1869 38913 1903 38947
rect 1903 38913 1912 38947
rect 1860 38904 1912 38913
rect 2780 38904 2832 38956
rect 2872 38904 2924 38956
rect 2412 38836 2464 38888
rect 4068 39040 4120 39092
rect 9864 39040 9916 39092
rect 3700 38972 3752 39024
rect 3792 38947 3844 38956
rect 3792 38913 3801 38947
rect 3801 38913 3835 38947
rect 3835 38913 3844 38947
rect 3792 38904 3844 38913
rect 3976 38904 4028 38956
rect 4068 38904 4120 38956
rect 4436 38947 4488 38956
rect 4436 38913 4445 38947
rect 4445 38913 4479 38947
rect 4479 38913 4488 38947
rect 4436 38904 4488 38913
rect 4988 38904 5040 38956
rect 1860 38768 1912 38820
rect 2780 38768 2832 38820
rect 3608 38768 3660 38820
rect 7012 38700 7064 38752
rect 10048 38743 10100 38752
rect 10048 38709 10057 38743
rect 10057 38709 10091 38743
rect 10091 38709 10100 38743
rect 10048 38700 10100 38709
rect 2582 38598 2634 38650
rect 2646 38598 2698 38650
rect 2710 38598 2762 38650
rect 2774 38598 2826 38650
rect 2838 38598 2890 38650
rect 5845 38598 5897 38650
rect 5909 38598 5961 38650
rect 5973 38598 6025 38650
rect 6037 38598 6089 38650
rect 6101 38598 6153 38650
rect 9109 38598 9161 38650
rect 9173 38598 9225 38650
rect 9237 38598 9289 38650
rect 9301 38598 9353 38650
rect 9365 38598 9417 38650
rect 2780 38292 2832 38344
rect 3240 38496 3292 38548
rect 3516 38428 3568 38480
rect 3240 38360 3292 38412
rect 3516 38292 3568 38344
rect 4344 38360 4396 38412
rect 4436 38292 4488 38344
rect 4988 38224 5040 38276
rect 2136 38199 2188 38208
rect 2136 38165 2145 38199
rect 2145 38165 2179 38199
rect 2179 38165 2188 38199
rect 2136 38156 2188 38165
rect 2228 38156 2280 38208
rect 4068 38156 4120 38208
rect 4213 38054 4265 38106
rect 4277 38054 4329 38106
rect 4341 38054 4393 38106
rect 4405 38054 4457 38106
rect 4469 38054 4521 38106
rect 7477 38054 7529 38106
rect 7541 38054 7593 38106
rect 7605 38054 7657 38106
rect 7669 38054 7721 38106
rect 7733 38054 7785 38106
rect 1768 37952 1820 38004
rect 5632 37884 5684 37936
rect 2780 37816 2832 37868
rect 9864 37859 9916 37868
rect 9864 37825 9873 37859
rect 9873 37825 9907 37859
rect 9907 37825 9916 37859
rect 9864 37816 9916 37825
rect 2228 37680 2280 37732
rect 7288 37680 7340 37732
rect 1492 37655 1544 37664
rect 1492 37621 1501 37655
rect 1501 37621 1535 37655
rect 1535 37621 1544 37655
rect 1492 37612 1544 37621
rect 10048 37655 10100 37664
rect 10048 37621 10057 37655
rect 10057 37621 10091 37655
rect 10091 37621 10100 37655
rect 10048 37612 10100 37621
rect 2582 37510 2634 37562
rect 2646 37510 2698 37562
rect 2710 37510 2762 37562
rect 2774 37510 2826 37562
rect 2838 37510 2890 37562
rect 5845 37510 5897 37562
rect 5909 37510 5961 37562
rect 5973 37510 6025 37562
rect 6037 37510 6089 37562
rect 6101 37510 6153 37562
rect 9109 37510 9161 37562
rect 9173 37510 9225 37562
rect 9237 37510 9289 37562
rect 9301 37510 9353 37562
rect 9365 37510 9417 37562
rect 2320 37451 2372 37460
rect 2320 37417 2329 37451
rect 2329 37417 2363 37451
rect 2363 37417 2372 37451
rect 2320 37408 2372 37417
rect 2136 37340 2188 37392
rect 1584 37204 1636 37256
rect 2320 37272 2372 37324
rect 2136 37204 2188 37256
rect 3424 37204 3476 37256
rect 3976 37204 4028 37256
rect 1676 37111 1728 37120
rect 1676 37077 1685 37111
rect 1685 37077 1719 37111
rect 1719 37077 1728 37111
rect 1676 37068 1728 37077
rect 2780 37068 2832 37120
rect 8760 37068 8812 37120
rect 10048 37111 10100 37120
rect 10048 37077 10057 37111
rect 10057 37077 10091 37111
rect 10091 37077 10100 37111
rect 10048 37068 10100 37077
rect 4213 36966 4265 37018
rect 4277 36966 4329 37018
rect 4341 36966 4393 37018
rect 4405 36966 4457 37018
rect 4469 36966 4521 37018
rect 7477 36966 7529 37018
rect 7541 36966 7593 37018
rect 7605 36966 7657 37018
rect 7669 36966 7721 37018
rect 7733 36966 7785 37018
rect 1676 36864 1728 36916
rect 9864 36864 9916 36916
rect 5540 36796 5592 36848
rect 2228 36728 2280 36780
rect 2780 36728 2832 36780
rect 3516 36728 3568 36780
rect 3792 36771 3844 36780
rect 3792 36737 3801 36771
rect 3801 36737 3835 36771
rect 3835 36737 3844 36771
rect 3792 36728 3844 36737
rect 3056 36635 3108 36644
rect 3056 36601 3065 36635
rect 3065 36601 3099 36635
rect 3099 36601 3108 36635
rect 3056 36592 3108 36601
rect 4896 36660 4948 36712
rect 5448 36660 5500 36712
rect 204 36524 256 36576
rect 940 36524 992 36576
rect 1400 36524 1452 36576
rect 2228 36567 2280 36576
rect 2228 36533 2237 36567
rect 2237 36533 2271 36567
rect 2271 36533 2280 36567
rect 2228 36524 2280 36533
rect 5080 36524 5132 36576
rect 5448 36524 5500 36576
rect 7932 36524 7984 36576
rect 8116 36524 8168 36576
rect 2582 36422 2634 36474
rect 2646 36422 2698 36474
rect 2710 36422 2762 36474
rect 2774 36422 2826 36474
rect 2838 36422 2890 36474
rect 5845 36422 5897 36474
rect 5909 36422 5961 36474
rect 5973 36422 6025 36474
rect 6037 36422 6089 36474
rect 6101 36422 6153 36474
rect 9109 36422 9161 36474
rect 9173 36422 9225 36474
rect 9237 36422 9289 36474
rect 9301 36422 9353 36474
rect 9365 36422 9417 36474
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 5172 36320 5224 36372
rect 5540 36320 5592 36372
rect 3424 36252 3476 36304
rect 3792 36252 3844 36304
rect 8576 36184 8628 36236
rect 3516 36116 3568 36168
rect 3884 36116 3936 36168
rect 9864 36159 9916 36168
rect 9864 36125 9873 36159
rect 9873 36125 9907 36159
rect 9907 36125 9916 36159
rect 9864 36116 9916 36125
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 10048 36023 10100 36032
rect 10048 35989 10057 36023
rect 10057 35989 10091 36023
rect 10091 35989 10100 36023
rect 10048 35980 10100 35989
rect 4213 35878 4265 35930
rect 4277 35878 4329 35930
rect 4341 35878 4393 35930
rect 4405 35878 4457 35930
rect 4469 35878 4521 35930
rect 7477 35878 7529 35930
rect 7541 35878 7593 35930
rect 7605 35878 7657 35930
rect 7669 35878 7721 35930
rect 7733 35878 7785 35930
rect 6920 35776 6972 35828
rect 2320 35708 2372 35760
rect 1768 35683 1820 35692
rect 1768 35649 1777 35683
rect 1777 35649 1811 35683
rect 1811 35649 1820 35683
rect 1768 35640 1820 35649
rect 2412 35640 2464 35692
rect 3516 35708 3568 35760
rect 3608 35640 3660 35692
rect 9772 35640 9824 35692
rect 4160 35572 4212 35624
rect 8852 35504 8904 35556
rect 4988 35436 5040 35488
rect 5356 35436 5408 35488
rect 10048 35479 10100 35488
rect 10048 35445 10057 35479
rect 10057 35445 10091 35479
rect 10091 35445 10100 35479
rect 10048 35436 10100 35445
rect 2582 35334 2634 35386
rect 2646 35334 2698 35386
rect 2710 35334 2762 35386
rect 2774 35334 2826 35386
rect 2838 35334 2890 35386
rect 5845 35334 5897 35386
rect 5909 35334 5961 35386
rect 5973 35334 6025 35386
rect 6037 35334 6089 35386
rect 6101 35334 6153 35386
rect 9109 35334 9161 35386
rect 9173 35334 9225 35386
rect 9237 35334 9289 35386
rect 9301 35334 9353 35386
rect 9365 35334 9417 35386
rect 9772 35232 9824 35284
rect 8392 35164 8444 35216
rect 6276 35096 6328 35148
rect 2412 35071 2464 35080
rect 2412 35037 2421 35071
rect 2421 35037 2455 35071
rect 2455 35037 2464 35071
rect 2412 35028 2464 35037
rect 3424 35028 3476 35080
rect 4160 35028 4212 35080
rect 9772 35028 9824 35080
rect 1492 34935 1544 34944
rect 1492 34901 1501 34935
rect 1501 34901 1535 34935
rect 1535 34901 1544 34935
rect 1492 34892 1544 34901
rect 10048 34935 10100 34944
rect 10048 34901 10057 34935
rect 10057 34901 10091 34935
rect 10091 34901 10100 34935
rect 10048 34892 10100 34901
rect 4213 34790 4265 34842
rect 4277 34790 4329 34842
rect 4341 34790 4393 34842
rect 4405 34790 4457 34842
rect 4469 34790 4521 34842
rect 7477 34790 7529 34842
rect 7541 34790 7593 34842
rect 7605 34790 7657 34842
rect 7669 34790 7721 34842
rect 7733 34790 7785 34842
rect 1584 34688 1636 34740
rect 8668 34620 8720 34672
rect 1584 34595 1636 34604
rect 1584 34561 1593 34595
rect 1593 34561 1627 34595
rect 1627 34561 1636 34595
rect 1584 34552 1636 34561
rect 2228 34595 2280 34604
rect 2228 34561 2237 34595
rect 2237 34561 2271 34595
rect 2271 34561 2280 34595
rect 2228 34552 2280 34561
rect 2412 34595 2464 34604
rect 2412 34561 2421 34595
rect 2421 34561 2455 34595
rect 2455 34561 2464 34595
rect 2412 34552 2464 34561
rect 3240 34552 3292 34604
rect 3240 34391 3292 34400
rect 3240 34357 3249 34391
rect 3249 34357 3283 34391
rect 3283 34357 3292 34391
rect 3240 34348 3292 34357
rect 2582 34246 2634 34298
rect 2646 34246 2698 34298
rect 2710 34246 2762 34298
rect 2774 34246 2826 34298
rect 2838 34246 2890 34298
rect 5845 34246 5897 34298
rect 5909 34246 5961 34298
rect 5973 34246 6025 34298
rect 6037 34246 6089 34298
rect 6101 34246 6153 34298
rect 9109 34246 9161 34298
rect 9173 34246 9225 34298
rect 9237 34246 9289 34298
rect 9301 34246 9353 34298
rect 9365 34246 9417 34298
rect 1768 34144 1820 34196
rect 2228 34144 2280 34196
rect 9864 34144 9916 34196
rect 3056 34119 3108 34128
rect 3056 34085 3065 34119
rect 3065 34085 3099 34119
rect 3099 34085 3108 34119
rect 3056 34076 3108 34085
rect 1952 33940 2004 33992
rect 3332 33940 3384 33992
rect 3424 33872 3476 33924
rect 9680 33940 9732 33992
rect 1492 33847 1544 33856
rect 1492 33813 1501 33847
rect 1501 33813 1535 33847
rect 1535 33813 1544 33847
rect 1492 33804 1544 33813
rect 2320 33847 2372 33856
rect 2320 33813 2329 33847
rect 2329 33813 2363 33847
rect 2363 33813 2372 33847
rect 2320 33804 2372 33813
rect 5356 33804 5408 33856
rect 5540 33804 5592 33856
rect 10048 33847 10100 33856
rect 10048 33813 10057 33847
rect 10057 33813 10091 33847
rect 10091 33813 10100 33847
rect 10048 33804 10100 33813
rect 4213 33702 4265 33754
rect 4277 33702 4329 33754
rect 4341 33702 4393 33754
rect 4405 33702 4457 33754
rect 4469 33702 4521 33754
rect 7477 33702 7529 33754
rect 7541 33702 7593 33754
rect 7605 33702 7657 33754
rect 7669 33702 7721 33754
rect 7733 33702 7785 33754
rect 9772 33600 9824 33652
rect 1952 33464 2004 33516
rect 2412 33464 2464 33516
rect 2504 33464 2556 33516
rect 2228 33396 2280 33448
rect 3424 33464 3476 33516
rect 7104 33464 7156 33516
rect 9864 33507 9916 33516
rect 9864 33473 9873 33507
rect 9873 33473 9907 33507
rect 9907 33473 9916 33507
rect 9864 33464 9916 33473
rect 1400 33260 1452 33312
rect 10048 33303 10100 33312
rect 10048 33269 10057 33303
rect 10057 33269 10091 33303
rect 10091 33269 10100 33303
rect 10048 33260 10100 33269
rect 2582 33158 2634 33210
rect 2646 33158 2698 33210
rect 2710 33158 2762 33210
rect 2774 33158 2826 33210
rect 2838 33158 2890 33210
rect 5845 33158 5897 33210
rect 5909 33158 5961 33210
rect 5973 33158 6025 33210
rect 6037 33158 6089 33210
rect 6101 33158 6153 33210
rect 9109 33158 9161 33210
rect 9173 33158 9225 33210
rect 9237 33158 9289 33210
rect 9301 33158 9353 33210
rect 9365 33158 9417 33210
rect 2964 33056 3016 33108
rect 4804 33056 4856 33108
rect 2320 32920 2372 32972
rect 2504 32920 2556 32972
rect 1216 32852 1268 32904
rect 2044 32852 2096 32904
rect 4804 32920 4856 32972
rect 5540 32852 5592 32904
rect 1216 32716 1268 32768
rect 2320 32759 2372 32768
rect 2320 32725 2329 32759
rect 2329 32725 2363 32759
rect 2363 32725 2372 32759
rect 2320 32716 2372 32725
rect 4213 32614 4265 32666
rect 4277 32614 4329 32666
rect 4341 32614 4393 32666
rect 4405 32614 4457 32666
rect 4469 32614 4521 32666
rect 7477 32614 7529 32666
rect 7541 32614 7593 32666
rect 7605 32614 7657 32666
rect 7669 32614 7721 32666
rect 7733 32614 7785 32666
rect 1308 32512 1360 32564
rect 1308 32376 1360 32428
rect 2504 32512 2556 32564
rect 9680 32512 9732 32564
rect 1952 32444 2004 32496
rect 2136 32419 2188 32428
rect 2136 32385 2145 32419
rect 2145 32385 2179 32419
rect 2179 32385 2188 32419
rect 2136 32376 2188 32385
rect 6552 32444 6604 32496
rect 3424 32419 3476 32428
rect 3424 32385 3433 32419
rect 3433 32385 3467 32419
rect 3467 32385 3476 32419
rect 3424 32376 3476 32385
rect 3976 32376 4028 32428
rect 10048 32283 10100 32292
rect 10048 32249 10057 32283
rect 10057 32249 10091 32283
rect 10091 32249 10100 32283
rect 10048 32240 10100 32249
rect 1492 32172 1544 32224
rect 2320 32172 2372 32224
rect 2582 32070 2634 32122
rect 2646 32070 2698 32122
rect 2710 32070 2762 32122
rect 2774 32070 2826 32122
rect 2838 32070 2890 32122
rect 5845 32070 5897 32122
rect 5909 32070 5961 32122
rect 5973 32070 6025 32122
rect 6037 32070 6089 32122
rect 6101 32070 6153 32122
rect 9109 32070 9161 32122
rect 9173 32070 9225 32122
rect 9237 32070 9289 32122
rect 9301 32070 9353 32122
rect 9365 32070 9417 32122
rect 1492 31968 1544 32020
rect 9864 31968 9916 32020
rect 2320 31832 2372 31884
rect 3424 31764 3476 31816
rect 3976 31807 4028 31816
rect 3976 31773 3985 31807
rect 3985 31773 4019 31807
rect 4019 31773 4028 31807
rect 3976 31764 4028 31773
rect 4068 31764 4120 31816
rect 7196 31764 7248 31816
rect 3608 31696 3660 31748
rect 2412 31671 2464 31680
rect 2412 31637 2421 31671
rect 2421 31637 2455 31671
rect 2455 31637 2464 31671
rect 2412 31628 2464 31637
rect 3976 31628 4028 31680
rect 10048 31671 10100 31680
rect 10048 31637 10057 31671
rect 10057 31637 10091 31671
rect 10091 31637 10100 31671
rect 10048 31628 10100 31637
rect 4213 31526 4265 31578
rect 4277 31526 4329 31578
rect 4341 31526 4393 31578
rect 4405 31526 4457 31578
rect 4469 31526 4521 31578
rect 7477 31526 7529 31578
rect 7541 31526 7593 31578
rect 7605 31526 7657 31578
rect 7669 31526 7721 31578
rect 7733 31526 7785 31578
rect 940 31356 992 31408
rect 3056 31220 3108 31272
rect 2412 31127 2464 31136
rect 2412 31093 2421 31127
rect 2421 31093 2455 31127
rect 2455 31093 2464 31127
rect 2412 31084 2464 31093
rect 10048 31127 10100 31136
rect 10048 31093 10057 31127
rect 10057 31093 10091 31127
rect 10091 31093 10100 31127
rect 10048 31084 10100 31093
rect 2582 30982 2634 31034
rect 2646 30982 2698 31034
rect 2710 30982 2762 31034
rect 2774 30982 2826 31034
rect 2838 30982 2890 31034
rect 5845 30982 5897 31034
rect 5909 30982 5961 31034
rect 5973 30982 6025 31034
rect 6037 30982 6089 31034
rect 6101 30982 6153 31034
rect 9109 30982 9161 31034
rect 9173 30982 9225 31034
rect 9237 30982 9289 31034
rect 9301 30982 9353 31034
rect 9365 30982 9417 31034
rect 296 30676 348 30728
rect 2320 30719 2372 30728
rect 2320 30685 2329 30719
rect 2329 30685 2363 30719
rect 2363 30685 2372 30719
rect 2320 30676 2372 30685
rect 1492 30583 1544 30592
rect 1492 30549 1501 30583
rect 1501 30549 1535 30583
rect 1535 30549 1544 30583
rect 1492 30540 1544 30549
rect 1768 30540 1820 30592
rect 4213 30438 4265 30490
rect 4277 30438 4329 30490
rect 4341 30438 4393 30490
rect 4405 30438 4457 30490
rect 4469 30438 4521 30490
rect 7477 30438 7529 30490
rect 7541 30438 7593 30490
rect 7605 30438 7657 30490
rect 7669 30438 7721 30490
rect 7733 30438 7785 30490
rect 1492 30336 1544 30388
rect 1676 30336 1728 30388
rect 1860 30268 1912 30320
rect 1676 30243 1728 30252
rect 1676 30209 1685 30243
rect 1685 30209 1719 30243
rect 1719 30209 1728 30243
rect 1676 30200 1728 30209
rect 1860 30132 1912 30184
rect 2136 30336 2188 30388
rect 2136 30243 2188 30252
rect 2136 30209 2145 30243
rect 2145 30209 2179 30243
rect 2179 30209 2188 30243
rect 2136 30200 2188 30209
rect 2964 30243 3016 30252
rect 2964 30209 2973 30243
rect 2973 30209 3007 30243
rect 3007 30209 3016 30243
rect 2964 30200 3016 30209
rect 9864 30243 9916 30252
rect 9864 30209 9873 30243
rect 9873 30209 9907 30243
rect 9907 30209 9916 30243
rect 9864 30200 9916 30209
rect 2044 30064 2096 30116
rect 1400 29996 1452 30048
rect 10048 30039 10100 30048
rect 10048 30005 10057 30039
rect 10057 30005 10091 30039
rect 10091 30005 10100 30039
rect 10048 29996 10100 30005
rect 2582 29894 2634 29946
rect 2646 29894 2698 29946
rect 2710 29894 2762 29946
rect 2774 29894 2826 29946
rect 2838 29894 2890 29946
rect 5845 29894 5897 29946
rect 5909 29894 5961 29946
rect 5973 29894 6025 29946
rect 6037 29894 6089 29946
rect 6101 29894 6153 29946
rect 9109 29894 9161 29946
rect 9173 29894 9225 29946
rect 9237 29894 9289 29946
rect 9301 29894 9353 29946
rect 9365 29894 9417 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 1676 29792 1728 29844
rect 3056 29792 3108 29844
rect 1584 29656 1636 29708
rect 1768 29631 1820 29640
rect 1768 29597 1777 29631
rect 1777 29597 1811 29631
rect 1811 29597 1820 29631
rect 1768 29588 1820 29597
rect 2964 29588 3016 29640
rect 3056 29631 3108 29640
rect 3056 29597 3065 29631
rect 3065 29597 3099 29631
rect 3099 29597 3108 29631
rect 3056 29588 3108 29597
rect 3240 29452 3292 29504
rect 3700 29452 3752 29504
rect 4213 29350 4265 29402
rect 4277 29350 4329 29402
rect 4341 29350 4393 29402
rect 4405 29350 4457 29402
rect 4469 29350 4521 29402
rect 7477 29350 7529 29402
rect 7541 29350 7593 29402
rect 7605 29350 7657 29402
rect 7669 29350 7721 29402
rect 7733 29350 7785 29402
rect 2044 29248 2096 29300
rect 2412 29248 2464 29300
rect 2780 29180 2832 29232
rect 2412 29112 2464 29164
rect 3424 29248 3476 29300
rect 10968 29223 11020 29232
rect 10968 29189 10977 29223
rect 10977 29189 11011 29223
rect 11011 29189 11020 29223
rect 10968 29180 11020 29189
rect 3792 29155 3844 29164
rect 3792 29121 3801 29155
rect 3801 29121 3835 29155
rect 3835 29121 3844 29155
rect 3792 29112 3844 29121
rect 8024 29044 8076 29096
rect 4068 28976 4120 29028
rect 1400 28908 1452 28960
rect 2964 28908 3016 28960
rect 3056 28908 3108 28960
rect 3424 28908 3476 28960
rect 4896 28908 4948 28960
rect 5080 28908 5132 28960
rect 10140 28951 10192 28960
rect 10140 28917 10149 28951
rect 10149 28917 10183 28951
rect 10183 28917 10192 28951
rect 10140 28908 10192 28917
rect 2582 28806 2634 28858
rect 2646 28806 2698 28858
rect 2710 28806 2762 28858
rect 2774 28806 2826 28858
rect 2838 28806 2890 28858
rect 5845 28806 5897 28858
rect 5909 28806 5961 28858
rect 5973 28806 6025 28858
rect 6037 28806 6089 28858
rect 6101 28806 6153 28858
rect 9109 28806 9161 28858
rect 9173 28806 9225 28858
rect 9237 28806 9289 28858
rect 9301 28806 9353 28858
rect 9365 28806 9417 28858
rect 388 28704 440 28756
rect 4620 28704 4672 28756
rect 4896 28704 4948 28756
rect 5448 28636 5500 28688
rect 2780 28543 2832 28552
rect 2780 28509 2789 28543
rect 2789 28509 2823 28543
rect 2823 28509 2832 28543
rect 3976 28543 4028 28552
rect 2780 28500 2832 28509
rect 3976 28509 3985 28543
rect 3985 28509 4019 28543
rect 4019 28509 4028 28543
rect 3976 28500 4028 28509
rect 4712 28432 4764 28484
rect 2688 28364 2740 28416
rect 4213 28262 4265 28314
rect 4277 28262 4329 28314
rect 4341 28262 4393 28314
rect 4405 28262 4457 28314
rect 4469 28262 4521 28314
rect 7477 28262 7529 28314
rect 7541 28262 7593 28314
rect 7605 28262 7657 28314
rect 7669 28262 7721 28314
rect 7733 28262 7785 28314
rect 2780 28160 2832 28212
rect 1492 28135 1544 28144
rect 1492 28101 1501 28135
rect 1501 28101 1535 28135
rect 1535 28101 1544 28135
rect 1492 28092 1544 28101
rect 2688 28092 2740 28144
rect 2320 28067 2372 28076
rect 2320 28033 2329 28067
rect 2329 28033 2363 28067
rect 2363 28033 2372 28067
rect 2320 28024 2372 28033
rect 2412 28024 2464 28076
rect 3056 28024 3108 28076
rect 3424 28024 3476 28076
rect 4620 27888 4672 27940
rect 1952 27820 2004 27872
rect 2582 27718 2634 27770
rect 2646 27718 2698 27770
rect 2710 27718 2762 27770
rect 2774 27718 2826 27770
rect 2838 27718 2890 27770
rect 5845 27718 5897 27770
rect 5909 27718 5961 27770
rect 5973 27718 6025 27770
rect 6037 27718 6089 27770
rect 6101 27718 6153 27770
rect 9109 27718 9161 27770
rect 9173 27718 9225 27770
rect 9237 27718 9289 27770
rect 9301 27718 9353 27770
rect 9365 27718 9417 27770
rect 2412 27616 2464 27668
rect 3792 27616 3844 27668
rect 10140 27616 10192 27668
rect 2872 27480 2924 27532
rect 9864 27548 9916 27600
rect 7380 27480 7432 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 2136 27455 2188 27464
rect 2136 27421 2145 27455
rect 2145 27421 2179 27455
rect 2179 27421 2188 27455
rect 2136 27412 2188 27421
rect 2320 27455 2372 27464
rect 2320 27421 2329 27455
rect 2329 27421 2363 27455
rect 2363 27421 2372 27455
rect 2320 27412 2372 27421
rect 2596 27412 2648 27464
rect 2780 27344 2832 27396
rect 3792 27455 3844 27464
rect 3792 27421 3807 27455
rect 3807 27421 3841 27455
rect 3841 27421 3844 27455
rect 3792 27412 3844 27421
rect 3976 27455 4028 27464
rect 3976 27421 3985 27455
rect 3985 27421 4019 27455
rect 4019 27421 4028 27455
rect 3976 27412 4028 27421
rect 4620 27412 4672 27464
rect 6276 27344 6328 27396
rect 1860 27276 1912 27328
rect 2872 27276 2924 27328
rect 5724 27276 5776 27328
rect 4213 27174 4265 27226
rect 4277 27174 4329 27226
rect 4341 27174 4393 27226
rect 4405 27174 4457 27226
rect 4469 27174 4521 27226
rect 7477 27174 7529 27226
rect 7541 27174 7593 27226
rect 7605 27174 7657 27226
rect 7669 27174 7721 27226
rect 7733 27174 7785 27226
rect 2320 27072 2372 27124
rect 664 27004 716 27056
rect 3516 27072 3568 27124
rect 4068 27072 4120 27124
rect 4712 27072 4764 27124
rect 1952 26936 2004 26988
rect 2596 26979 2648 26988
rect 2596 26945 2605 26979
rect 2605 26945 2639 26979
rect 2639 26945 2648 26979
rect 2596 26936 2648 26945
rect 3056 26936 3108 26988
rect 2228 26868 2280 26920
rect 2872 26800 2924 26852
rect 4620 26936 4672 26988
rect 10140 26979 10192 26988
rect 3700 26868 3752 26920
rect 10140 26945 10149 26979
rect 10149 26945 10183 26979
rect 10183 26945 10192 26979
rect 10140 26936 10192 26945
rect 3608 26732 3660 26784
rect 2582 26630 2634 26682
rect 2646 26630 2698 26682
rect 2710 26630 2762 26682
rect 2774 26630 2826 26682
rect 2838 26630 2890 26682
rect 5845 26630 5897 26682
rect 5909 26630 5961 26682
rect 5973 26630 6025 26682
rect 6037 26630 6089 26682
rect 6101 26630 6153 26682
rect 9109 26630 9161 26682
rect 9173 26630 9225 26682
rect 9237 26630 9289 26682
rect 9301 26630 9353 26682
rect 9365 26630 9417 26682
rect 1952 26528 2004 26580
rect 2412 26460 2464 26512
rect 2596 26460 2648 26512
rect 1584 26392 1636 26444
rect 1952 26392 2004 26444
rect 1216 26324 1268 26376
rect 1492 26324 1544 26376
rect 2136 26324 2188 26376
rect 3516 26324 3568 26376
rect 4712 26256 4764 26308
rect 1584 26231 1636 26240
rect 1584 26197 1593 26231
rect 1593 26197 1627 26231
rect 1627 26197 1636 26231
rect 1584 26188 1636 26197
rect 2320 26188 2372 26240
rect 4213 26086 4265 26138
rect 4277 26086 4329 26138
rect 4341 26086 4393 26138
rect 4405 26086 4457 26138
rect 4469 26086 4521 26138
rect 7477 26086 7529 26138
rect 7541 26086 7593 26138
rect 7605 26086 7657 26138
rect 7669 26086 7721 26138
rect 7733 26086 7785 26138
rect 4896 25916 4948 25968
rect 1860 25891 1912 25900
rect 1860 25857 1869 25891
rect 1869 25857 1903 25891
rect 1903 25857 1912 25891
rect 1860 25848 1912 25857
rect 2964 25848 3016 25900
rect 2596 25780 2648 25832
rect 1860 25712 1912 25764
rect 2044 25644 2096 25696
rect 2582 25542 2634 25594
rect 2646 25542 2698 25594
rect 2710 25542 2762 25594
rect 2774 25542 2826 25594
rect 2838 25542 2890 25594
rect 5845 25542 5897 25594
rect 5909 25542 5961 25594
rect 5973 25542 6025 25594
rect 6037 25542 6089 25594
rect 6101 25542 6153 25594
rect 9109 25542 9161 25594
rect 9173 25542 9225 25594
rect 9237 25542 9289 25594
rect 9301 25542 9353 25594
rect 9365 25542 9417 25594
rect 1124 25440 1176 25492
rect 4988 25440 5040 25492
rect 10140 25483 10192 25492
rect 10140 25449 10149 25483
rect 10149 25449 10183 25483
rect 10183 25449 10192 25483
rect 10140 25440 10192 25449
rect 3240 25372 3292 25424
rect 3516 25372 3568 25424
rect 2044 25236 2096 25288
rect 2320 25279 2372 25288
rect 2320 25245 2329 25279
rect 2329 25245 2363 25279
rect 2363 25245 2372 25279
rect 2320 25236 2372 25245
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 2872 25100 2924 25152
rect 4213 24998 4265 25050
rect 4277 24998 4329 25050
rect 4341 24998 4393 25050
rect 4405 24998 4457 25050
rect 4469 24998 4521 25050
rect 7477 24998 7529 25050
rect 7541 24998 7593 25050
rect 7605 24998 7657 25050
rect 7669 24998 7721 25050
rect 7733 24998 7785 25050
rect 2320 24896 2372 24948
rect 2596 24896 2648 24948
rect 3332 24828 3384 24880
rect 10232 24828 10284 24880
rect 1492 24760 1544 24812
rect 2872 24760 2924 24812
rect 572 24692 624 24744
rect 4620 24760 4672 24812
rect 2964 24624 3016 24676
rect 5172 24624 5224 24676
rect 2582 24454 2634 24506
rect 2646 24454 2698 24506
rect 2710 24454 2762 24506
rect 2774 24454 2826 24506
rect 2838 24454 2890 24506
rect 5845 24454 5897 24506
rect 5909 24454 5961 24506
rect 5973 24454 6025 24506
rect 6037 24454 6089 24506
rect 6101 24454 6153 24506
rect 9109 24454 9161 24506
rect 9173 24454 9225 24506
rect 9237 24454 9289 24506
rect 9301 24454 9353 24506
rect 9365 24454 9417 24506
rect 5080 24352 5132 24404
rect 10140 24395 10192 24404
rect 10140 24361 10149 24395
rect 10149 24361 10183 24395
rect 10183 24361 10192 24395
rect 10140 24352 10192 24361
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 1584 24148 1636 24200
rect 3148 24191 3200 24200
rect 3148 24157 3157 24191
rect 3157 24157 3191 24191
rect 3191 24157 3200 24191
rect 3148 24148 3200 24157
rect 2136 24012 2188 24064
rect 2504 24012 2556 24064
rect 4213 23910 4265 23962
rect 4277 23910 4329 23962
rect 4341 23910 4393 23962
rect 4405 23910 4457 23962
rect 4469 23910 4521 23962
rect 7477 23910 7529 23962
rect 7541 23910 7593 23962
rect 7605 23910 7657 23962
rect 7669 23910 7721 23962
rect 7733 23910 7785 23962
rect 1032 23740 1084 23792
rect 1216 23672 1268 23724
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2504 23672 2556 23681
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 1584 23511 1636 23520
rect 1584 23477 1593 23511
rect 1593 23477 1627 23511
rect 1627 23477 1636 23511
rect 1584 23468 1636 23477
rect 10048 23511 10100 23520
rect 10048 23477 10057 23511
rect 10057 23477 10091 23511
rect 10091 23477 10100 23511
rect 10048 23468 10100 23477
rect 2582 23366 2634 23418
rect 2646 23366 2698 23418
rect 2710 23366 2762 23418
rect 2774 23366 2826 23418
rect 2838 23366 2890 23418
rect 5845 23366 5897 23418
rect 5909 23366 5961 23418
rect 5973 23366 6025 23418
rect 6037 23366 6089 23418
rect 6101 23366 6153 23418
rect 9109 23366 9161 23418
rect 9173 23366 9225 23418
rect 9237 23366 9289 23418
rect 9301 23366 9353 23418
rect 9365 23366 9417 23418
rect 2504 23264 2556 23316
rect 3792 23264 3844 23316
rect 9864 23264 9916 23316
rect 10140 23307 10192 23316
rect 10140 23273 10149 23307
rect 10149 23273 10183 23307
rect 10183 23273 10192 23307
rect 10140 23264 10192 23273
rect 3516 23196 3568 23248
rect 1584 23103 1636 23112
rect 1584 23069 1593 23103
rect 1593 23069 1627 23103
rect 1627 23069 1636 23103
rect 1584 23060 1636 23069
rect 2136 23103 2188 23112
rect 2136 23069 2145 23103
rect 2145 23069 2179 23103
rect 2179 23069 2188 23103
rect 2136 23060 2188 23069
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 2964 23060 3016 23069
rect 3516 23060 3568 23112
rect 4213 22822 4265 22874
rect 4277 22822 4329 22874
rect 4341 22822 4393 22874
rect 4405 22822 4457 22874
rect 4469 22822 4521 22874
rect 7477 22822 7529 22874
rect 7541 22822 7593 22874
rect 7605 22822 7657 22874
rect 7669 22822 7721 22874
rect 7733 22822 7785 22874
rect 5356 22720 5408 22772
rect 3792 22652 3844 22704
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 9864 22627 9916 22636
rect 9864 22593 9873 22627
rect 9873 22593 9907 22627
rect 9907 22593 9916 22627
rect 9864 22584 9916 22593
rect 3976 22380 4028 22432
rect 10048 22423 10100 22432
rect 10048 22389 10057 22423
rect 10057 22389 10091 22423
rect 10091 22389 10100 22423
rect 10048 22380 10100 22389
rect 2582 22278 2634 22330
rect 2646 22278 2698 22330
rect 2710 22278 2762 22330
rect 2774 22278 2826 22330
rect 2838 22278 2890 22330
rect 5845 22278 5897 22330
rect 5909 22278 5961 22330
rect 5973 22278 6025 22330
rect 6037 22278 6089 22330
rect 6101 22278 6153 22330
rect 9109 22278 9161 22330
rect 9173 22278 9225 22330
rect 9237 22278 9289 22330
rect 9301 22278 9353 22330
rect 9365 22278 9417 22330
rect 3792 22219 3844 22228
rect 3792 22185 3801 22219
rect 3801 22185 3835 22219
rect 3835 22185 3844 22219
rect 3792 22176 3844 22185
rect 3424 22040 3476 22092
rect 2872 22015 2924 22024
rect 2872 21981 2881 22015
rect 2881 21981 2915 22015
rect 2915 21981 2924 22015
rect 2872 21972 2924 21981
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 9956 21972 10008 22024
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 4213 21734 4265 21786
rect 4277 21734 4329 21786
rect 4341 21734 4393 21786
rect 4405 21734 4457 21786
rect 4469 21734 4521 21786
rect 7477 21734 7529 21786
rect 7541 21734 7593 21786
rect 7605 21734 7657 21786
rect 7669 21734 7721 21786
rect 7733 21734 7785 21786
rect 1768 21632 1820 21684
rect 2136 21632 2188 21684
rect 2320 21632 2372 21684
rect 3332 21564 3384 21616
rect 2320 21496 2372 21548
rect 3884 21539 3936 21548
rect 1768 21428 1820 21480
rect 3884 21505 3893 21539
rect 3893 21505 3927 21539
rect 3927 21505 3936 21539
rect 3884 21496 3936 21505
rect 2504 21403 2556 21412
rect 2504 21369 2513 21403
rect 2513 21369 2547 21403
rect 2547 21369 2556 21403
rect 2504 21360 2556 21369
rect 3148 21292 3200 21344
rect 2582 21190 2634 21242
rect 2646 21190 2698 21242
rect 2710 21190 2762 21242
rect 2774 21190 2826 21242
rect 2838 21190 2890 21242
rect 5845 21190 5897 21242
rect 5909 21190 5961 21242
rect 5973 21190 6025 21242
rect 6037 21190 6089 21242
rect 6101 21190 6153 21242
rect 9109 21190 9161 21242
rect 9173 21190 9225 21242
rect 9237 21190 9289 21242
rect 9301 21190 9353 21242
rect 9365 21190 9417 21242
rect 1952 21131 2004 21140
rect 1952 21097 1961 21131
rect 1961 21097 1995 21131
rect 1995 21097 2004 21131
rect 1952 21088 2004 21097
rect 2320 21088 2372 21140
rect 2780 21020 2832 21072
rect 5264 21020 5316 21072
rect 3700 20884 3752 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 9772 20884 9824 20936
rect 2504 20859 2556 20868
rect 2504 20825 2513 20859
rect 2513 20825 2547 20859
rect 2547 20825 2556 20859
rect 2504 20816 2556 20825
rect 1768 20748 1820 20800
rect 1952 20748 2004 20800
rect 2964 20748 3016 20800
rect 3516 20748 3568 20800
rect 10048 20791 10100 20800
rect 10048 20757 10057 20791
rect 10057 20757 10091 20791
rect 10091 20757 10100 20791
rect 10048 20748 10100 20757
rect 4213 20646 4265 20698
rect 4277 20646 4329 20698
rect 4341 20646 4393 20698
rect 4405 20646 4457 20698
rect 4469 20646 4521 20698
rect 7477 20646 7529 20698
rect 7541 20646 7593 20698
rect 7605 20646 7657 20698
rect 7669 20646 7721 20698
rect 7733 20646 7785 20698
rect 1676 20544 1728 20596
rect 3056 20544 3108 20596
rect 3700 20544 3752 20596
rect 4068 20544 4120 20596
rect 9864 20544 9916 20596
rect 3516 20476 3568 20528
rect 2320 20408 2372 20460
rect 2780 20451 2832 20460
rect 2780 20417 2789 20451
rect 2789 20417 2823 20451
rect 2823 20417 2832 20451
rect 3424 20451 3476 20460
rect 2780 20408 2832 20417
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 4068 20451 4120 20460
rect 4068 20417 4077 20451
rect 4077 20417 4111 20451
rect 4111 20417 4120 20451
rect 4068 20408 4120 20417
rect 9864 20451 9916 20460
rect 3884 20340 3936 20392
rect 9864 20417 9873 20451
rect 9873 20417 9907 20451
rect 9907 20417 9916 20451
rect 9864 20408 9916 20417
rect 3240 20247 3292 20256
rect 3240 20213 3249 20247
rect 3249 20213 3283 20247
rect 3283 20213 3292 20247
rect 3240 20204 3292 20213
rect 10048 20247 10100 20256
rect 10048 20213 10057 20247
rect 10057 20213 10091 20247
rect 10091 20213 10100 20247
rect 10048 20204 10100 20213
rect 2582 20102 2634 20154
rect 2646 20102 2698 20154
rect 2710 20102 2762 20154
rect 2774 20102 2826 20154
rect 2838 20102 2890 20154
rect 5845 20102 5897 20154
rect 5909 20102 5961 20154
rect 5973 20102 6025 20154
rect 6037 20102 6089 20154
rect 6101 20102 6153 20154
rect 9109 20102 9161 20154
rect 9173 20102 9225 20154
rect 9237 20102 9289 20154
rect 9301 20102 9353 20154
rect 9365 20102 9417 20154
rect 2412 20000 2464 20052
rect 3516 20000 3568 20052
rect 3240 19864 3292 19916
rect 3148 19796 3200 19848
rect 4620 19728 4672 19780
rect 4712 19660 4764 19712
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 4213 19558 4265 19610
rect 4277 19558 4329 19610
rect 4341 19558 4393 19610
rect 4405 19558 4457 19610
rect 4469 19558 4521 19610
rect 7477 19558 7529 19610
rect 7541 19558 7593 19610
rect 7605 19558 7657 19610
rect 7669 19558 7721 19610
rect 7733 19558 7785 19610
rect 2228 19456 2280 19508
rect 2412 19456 2464 19508
rect 3056 19456 3108 19508
rect 9956 19499 10008 19508
rect 9956 19465 9965 19499
rect 9965 19465 9999 19499
rect 9999 19465 10008 19499
rect 9956 19456 10008 19465
rect 3424 19388 3476 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2412 19363 2464 19372
rect 2412 19329 2421 19363
rect 2421 19329 2455 19363
rect 2455 19329 2464 19363
rect 2412 19320 2464 19329
rect 3056 19363 3108 19372
rect 3056 19329 3065 19363
rect 3065 19329 3099 19363
rect 3099 19329 3108 19363
rect 3056 19320 3108 19329
rect 10140 19363 10192 19372
rect 10140 19329 10149 19363
rect 10149 19329 10183 19363
rect 10183 19329 10192 19363
rect 10140 19320 10192 19329
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2582 19014 2634 19066
rect 2646 19014 2698 19066
rect 2710 19014 2762 19066
rect 2774 19014 2826 19066
rect 2838 19014 2890 19066
rect 5845 19014 5897 19066
rect 5909 19014 5961 19066
rect 5973 19014 6025 19066
rect 6037 19014 6089 19066
rect 6101 19014 6153 19066
rect 9109 19014 9161 19066
rect 9173 19014 9225 19066
rect 9237 19014 9289 19066
rect 9301 19014 9353 19066
rect 9365 19014 9417 19066
rect 2044 18912 2096 18964
rect 9772 18912 9824 18964
rect 2780 18708 2832 18760
rect 3240 18751 3292 18760
rect 3240 18717 3249 18751
rect 3249 18717 3283 18751
rect 3283 18717 3292 18751
rect 3240 18708 3292 18717
rect 2320 18640 2372 18692
rect 9956 18708 10008 18760
rect 1952 18572 2004 18624
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 4213 18470 4265 18522
rect 4277 18470 4329 18522
rect 4341 18470 4393 18522
rect 4405 18470 4457 18522
rect 4469 18470 4521 18522
rect 7477 18470 7529 18522
rect 7541 18470 7593 18522
rect 7605 18470 7657 18522
rect 7669 18470 7721 18522
rect 7733 18470 7785 18522
rect 1860 18368 1912 18420
rect 2412 18368 2464 18420
rect 1952 18232 2004 18284
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 3056 18232 3108 18284
rect 9772 18232 9824 18284
rect 2136 18164 2188 18216
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 2582 17926 2634 17978
rect 2646 17926 2698 17978
rect 2710 17926 2762 17978
rect 2774 17926 2826 17978
rect 2838 17926 2890 17978
rect 5845 17926 5897 17978
rect 5909 17926 5961 17978
rect 5973 17926 6025 17978
rect 6037 17926 6089 17978
rect 6101 17926 6153 17978
rect 9109 17926 9161 17978
rect 9173 17926 9225 17978
rect 9237 17926 9289 17978
rect 9301 17926 9353 17978
rect 9365 17926 9417 17978
rect 3608 17824 3660 17876
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 2964 17688 3016 17740
rect 3516 17688 3568 17740
rect 1584 17620 1636 17672
rect 2136 17620 2188 17672
rect 2320 17620 2372 17672
rect 9680 17620 9732 17672
rect 1952 17484 2004 17536
rect 2596 17527 2648 17536
rect 2596 17493 2605 17527
rect 2605 17493 2639 17527
rect 2639 17493 2648 17527
rect 2596 17484 2648 17493
rect 3884 17552 3936 17604
rect 2964 17484 3016 17536
rect 4213 17382 4265 17434
rect 4277 17382 4329 17434
rect 4341 17382 4393 17434
rect 4405 17382 4457 17434
rect 4469 17382 4521 17434
rect 7477 17382 7529 17434
rect 7541 17382 7593 17434
rect 7605 17382 7657 17434
rect 7669 17382 7721 17434
rect 7733 17382 7785 17434
rect 2228 17280 2280 17332
rect 2596 17212 2648 17264
rect 10140 17212 10192 17264
rect 1216 17144 1268 17196
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 10048 17051 10100 17060
rect 10048 17017 10057 17051
rect 10057 17017 10091 17051
rect 10091 17017 10100 17051
rect 10048 17008 10100 17017
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 1768 16940 1820 16992
rect 2582 16838 2634 16890
rect 2646 16838 2698 16890
rect 2710 16838 2762 16890
rect 2774 16838 2826 16890
rect 2838 16838 2890 16890
rect 5845 16838 5897 16890
rect 5909 16838 5961 16890
rect 5973 16838 6025 16890
rect 6037 16838 6089 16890
rect 6101 16838 6153 16890
rect 9109 16838 9161 16890
rect 9173 16838 9225 16890
rect 9237 16838 9289 16890
rect 9301 16838 9353 16890
rect 9365 16838 9417 16890
rect 3148 16736 3200 16788
rect 2964 16643 3016 16652
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 1124 16532 1176 16584
rect 9864 16575 9916 16584
rect 2320 16464 2372 16516
rect 1400 16396 1452 16448
rect 2504 16396 2556 16448
rect 2964 16464 3016 16516
rect 3056 16507 3108 16516
rect 3056 16473 3065 16507
rect 3065 16473 3099 16507
rect 3099 16473 3108 16507
rect 3056 16464 3108 16473
rect 9864 16541 9873 16575
rect 9873 16541 9907 16575
rect 9907 16541 9916 16575
rect 9864 16532 9916 16541
rect 9772 16396 9824 16448
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 4213 16294 4265 16346
rect 4277 16294 4329 16346
rect 4341 16294 4393 16346
rect 4405 16294 4457 16346
rect 4469 16294 4521 16346
rect 7477 16294 7529 16346
rect 7541 16294 7593 16346
rect 7605 16294 7657 16346
rect 7669 16294 7721 16346
rect 7733 16294 7785 16346
rect 2044 16192 2096 16244
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 1860 16056 1912 16108
rect 3240 16099 3292 16108
rect 3240 16065 3249 16099
rect 3249 16065 3283 16099
rect 3283 16065 3292 16099
rect 3240 16056 3292 16065
rect 4988 16056 5040 16108
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 2044 15852 2096 15904
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 2582 15750 2634 15802
rect 2646 15750 2698 15802
rect 2710 15750 2762 15802
rect 2774 15750 2826 15802
rect 2838 15750 2890 15802
rect 5845 15750 5897 15802
rect 5909 15750 5961 15802
rect 5973 15750 6025 15802
rect 6037 15750 6089 15802
rect 6101 15750 6153 15802
rect 9109 15750 9161 15802
rect 9173 15750 9225 15802
rect 9237 15750 9289 15802
rect 9301 15750 9353 15802
rect 9365 15750 9417 15802
rect 1676 15648 1728 15700
rect 3056 15648 3108 15700
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 2044 15512 2096 15564
rect 2320 15512 2372 15564
rect 4068 15512 4120 15564
rect 9680 15512 9732 15564
rect 1584 15487 1636 15496
rect 1584 15453 1593 15487
rect 1593 15453 1627 15487
rect 1627 15453 1636 15487
rect 1584 15444 1636 15453
rect 1768 15444 1820 15496
rect 2412 15308 2464 15360
rect 2596 15351 2648 15360
rect 2596 15317 2605 15351
rect 2605 15317 2639 15351
rect 2639 15317 2648 15351
rect 2596 15308 2648 15317
rect 4988 15308 5040 15360
rect 4213 15206 4265 15258
rect 4277 15206 4329 15258
rect 4341 15206 4393 15258
rect 4405 15206 4457 15258
rect 4469 15206 4521 15258
rect 7477 15206 7529 15258
rect 7541 15206 7593 15258
rect 7605 15206 7657 15258
rect 7669 15206 7721 15258
rect 7733 15206 7785 15258
rect 1492 15104 1544 15156
rect 2780 15104 2832 15156
rect 3240 15104 3292 15156
rect 3424 15104 3476 15156
rect 3608 15104 3660 15156
rect 9036 15104 9088 15156
rect 9864 15104 9916 15156
rect 1400 14900 1452 14952
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 2136 14968 2188 15020
rect 3056 14968 3108 15020
rect 3240 14968 3292 15020
rect 7932 15036 7984 15088
rect 3608 14968 3660 15020
rect 3700 14900 3752 14952
rect 3516 14832 3568 14884
rect 3884 14764 3936 14816
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 2582 14662 2634 14714
rect 2646 14662 2698 14714
rect 2710 14662 2762 14714
rect 2774 14662 2826 14714
rect 2838 14662 2890 14714
rect 5845 14662 5897 14714
rect 5909 14662 5961 14714
rect 5973 14662 6025 14714
rect 6037 14662 6089 14714
rect 6101 14662 6153 14714
rect 9109 14662 9161 14714
rect 9173 14662 9225 14714
rect 9237 14662 9289 14714
rect 9301 14662 9353 14714
rect 9365 14662 9417 14714
rect 1860 14560 1912 14612
rect 3700 14492 3752 14544
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 4712 14424 4764 14476
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4160 14356 4212 14408
rect 8944 14220 8996 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 4213 14118 4265 14170
rect 4277 14118 4329 14170
rect 4341 14118 4393 14170
rect 4405 14118 4457 14170
rect 4469 14118 4521 14170
rect 7477 14118 7529 14170
rect 7541 14118 7593 14170
rect 7605 14118 7657 14170
rect 7669 14118 7721 14170
rect 7733 14118 7785 14170
rect 3056 14016 3108 14068
rect 9864 14016 9916 14068
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 2136 13880 2188 13932
rect 9772 13948 9824 14000
rect 3056 13880 3108 13932
rect 3332 13880 3384 13932
rect 3608 13880 3660 13932
rect 3792 13923 3844 13932
rect 3792 13889 3801 13923
rect 3801 13889 3835 13923
rect 3835 13889 3844 13923
rect 3792 13880 3844 13889
rect 4160 13880 4212 13932
rect 3424 13812 3476 13864
rect 3884 13812 3936 13864
rect 3148 13744 3200 13796
rect 3332 13744 3384 13796
rect 3424 13676 3476 13728
rect 4068 13676 4120 13728
rect 2582 13574 2634 13626
rect 2646 13574 2698 13626
rect 2710 13574 2762 13626
rect 2774 13574 2826 13626
rect 2838 13574 2890 13626
rect 5845 13574 5897 13626
rect 5909 13574 5961 13626
rect 5973 13574 6025 13626
rect 6037 13574 6089 13626
rect 6101 13574 6153 13626
rect 9109 13574 9161 13626
rect 9173 13574 9225 13626
rect 9237 13574 9289 13626
rect 9301 13574 9353 13626
rect 9365 13574 9417 13626
rect 2964 13472 3016 13524
rect 2780 13404 2832 13456
rect 3240 13404 3292 13456
rect 1952 13336 2004 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 3516 13336 3568 13388
rect 3148 13268 3200 13320
rect 4620 13268 4672 13320
rect 9956 13268 10008 13320
rect 3240 13200 3292 13252
rect 10048 13175 10100 13184
rect 10048 13141 10057 13175
rect 10057 13141 10091 13175
rect 10091 13141 10100 13175
rect 10048 13132 10100 13141
rect 4213 13030 4265 13082
rect 4277 13030 4329 13082
rect 4341 13030 4393 13082
rect 4405 13030 4457 13082
rect 4469 13030 4521 13082
rect 7477 13030 7529 13082
rect 7541 13030 7593 13082
rect 7605 13030 7657 13082
rect 7669 13030 7721 13082
rect 7733 13030 7785 13082
rect 2964 12860 3016 12912
rect 2044 12792 2096 12844
rect 3148 12792 3200 12844
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 1492 12724 1544 12776
rect 2780 12724 2832 12776
rect 2872 12724 2924 12776
rect 3148 12656 3200 12708
rect 3516 12656 3568 12708
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 2582 12486 2634 12538
rect 2646 12486 2698 12538
rect 2710 12486 2762 12538
rect 2774 12486 2826 12538
rect 2838 12486 2890 12538
rect 5845 12486 5897 12538
rect 5909 12486 5961 12538
rect 5973 12486 6025 12538
rect 6037 12486 6089 12538
rect 6101 12486 6153 12538
rect 9109 12486 9161 12538
rect 9173 12486 9225 12538
rect 9237 12486 9289 12538
rect 9301 12486 9353 12538
rect 9365 12486 9417 12538
rect 7840 12384 7892 12436
rect 3424 12248 3476 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 3884 12180 3936 12232
rect 9772 12180 9824 12232
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 4213 11942 4265 11994
rect 4277 11942 4329 11994
rect 4341 11942 4393 11994
rect 4405 11942 4457 11994
rect 4469 11942 4521 11994
rect 7477 11942 7529 11994
rect 7541 11942 7593 11994
rect 7605 11942 7657 11994
rect 7669 11942 7721 11994
rect 7733 11942 7785 11994
rect 6184 11840 6236 11892
rect 9956 11883 10008 11892
rect 9956 11849 9965 11883
rect 9965 11849 9999 11883
rect 9999 11849 10008 11883
rect 9956 11840 10008 11849
rect 2228 11704 2280 11756
rect 3332 11704 3384 11756
rect 10140 11747 10192 11756
rect 10140 11713 10149 11747
rect 10149 11713 10183 11747
rect 10183 11713 10192 11747
rect 10140 11704 10192 11713
rect 1308 11636 1360 11688
rect 2582 11398 2634 11450
rect 2646 11398 2698 11450
rect 2710 11398 2762 11450
rect 2774 11398 2826 11450
rect 2838 11398 2890 11450
rect 5845 11398 5897 11450
rect 5909 11398 5961 11450
rect 5973 11398 6025 11450
rect 6037 11398 6089 11450
rect 6101 11398 6153 11450
rect 9109 11398 9161 11450
rect 9173 11398 9225 11450
rect 9237 11398 9289 11450
rect 9301 11398 9353 11450
rect 9365 11398 9417 11450
rect 8208 11296 8260 11348
rect 1584 11228 1636 11280
rect 6736 11228 6788 11280
rect 2412 11160 2464 11212
rect 3516 11160 3568 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2872 11092 2924 11144
rect 3884 11092 3936 11144
rect 10048 10999 10100 11008
rect 10048 10965 10057 10999
rect 10057 10965 10091 10999
rect 10091 10965 10100 10999
rect 10048 10956 10100 10965
rect 4213 10854 4265 10906
rect 4277 10854 4329 10906
rect 4341 10854 4393 10906
rect 4405 10854 4457 10906
rect 4469 10854 4521 10906
rect 7477 10854 7529 10906
rect 7541 10854 7593 10906
rect 7605 10854 7657 10906
rect 7669 10854 7721 10906
rect 7733 10854 7785 10906
rect 1768 10616 1820 10668
rect 2872 10616 2924 10668
rect 3700 10616 3752 10668
rect 1308 10548 1360 10600
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 2582 10310 2634 10362
rect 2646 10310 2698 10362
rect 2710 10310 2762 10362
rect 2774 10310 2826 10362
rect 2838 10310 2890 10362
rect 5845 10310 5897 10362
rect 5909 10310 5961 10362
rect 5973 10310 6025 10362
rect 6037 10310 6089 10362
rect 6101 10310 6153 10362
rect 9109 10310 9161 10362
rect 9173 10310 9225 10362
rect 9237 10310 9289 10362
rect 9301 10310 9353 10362
rect 9365 10310 9417 10362
rect 6644 10208 6696 10260
rect 2964 10140 3016 10192
rect 3148 10140 3200 10192
rect 2780 10072 2832 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 3148 10004 3200 10056
rect 4213 9766 4265 9818
rect 4277 9766 4329 9818
rect 4341 9766 4393 9818
rect 4405 9766 4457 9818
rect 4469 9766 4521 9818
rect 7477 9766 7529 9818
rect 7541 9766 7593 9818
rect 7605 9766 7657 9818
rect 7669 9766 7721 9818
rect 7733 9766 7785 9818
rect 3516 9664 3568 9716
rect 1768 9528 1820 9580
rect 10140 9596 10192 9648
rect 4068 9528 4120 9580
rect 8392 9528 8444 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 2780 9460 2832 9512
rect 3976 9460 4028 9512
rect 3424 9392 3476 9444
rect 10048 9435 10100 9444
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 2582 9222 2634 9274
rect 2646 9222 2698 9274
rect 2710 9222 2762 9274
rect 2774 9222 2826 9274
rect 2838 9222 2890 9274
rect 5845 9222 5897 9274
rect 5909 9222 5961 9274
rect 5973 9222 6025 9274
rect 6037 9222 6089 9274
rect 6101 9222 6153 9274
rect 9109 9222 9161 9274
rect 9173 9222 9225 9274
rect 9237 9222 9289 9274
rect 9301 9222 9353 9274
rect 9365 9222 9417 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 3424 9120 3476 9172
rect 3792 9120 3844 9172
rect 3332 8916 3384 8968
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 4068 8916 4120 8968
rect 2964 8848 3016 8900
rect 8392 8848 8444 8900
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 9220 8780 9272 8832
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 4213 8678 4265 8730
rect 4277 8678 4329 8730
rect 4341 8678 4393 8730
rect 4405 8678 4457 8730
rect 4469 8678 4521 8730
rect 7477 8678 7529 8730
rect 7541 8678 7593 8730
rect 7605 8678 7657 8730
rect 7669 8678 7721 8730
rect 7733 8678 7785 8730
rect 4068 8576 4120 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 3148 8440 3200 8492
rect 3700 8440 3752 8492
rect 4068 8440 4120 8492
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 2582 8134 2634 8186
rect 2646 8134 2698 8186
rect 2710 8134 2762 8186
rect 2774 8134 2826 8186
rect 2838 8134 2890 8186
rect 5845 8134 5897 8186
rect 5909 8134 5961 8186
rect 5973 8134 6025 8186
rect 6037 8134 6089 8186
rect 6101 8134 6153 8186
rect 9109 8134 9161 8186
rect 9173 8134 9225 8186
rect 9237 8134 9289 8186
rect 9301 8134 9353 8186
rect 9365 8134 9417 8186
rect 1768 7896 1820 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 4804 7760 4856 7812
rect 9036 7692 9088 7744
rect 4213 7590 4265 7642
rect 4277 7590 4329 7642
rect 4341 7590 4393 7642
rect 4405 7590 4457 7642
rect 4469 7590 4521 7642
rect 7477 7590 7529 7642
rect 7541 7590 7593 7642
rect 7605 7590 7657 7642
rect 7669 7590 7721 7642
rect 7733 7590 7785 7642
rect 3608 7488 3660 7540
rect 3240 7420 3292 7472
rect 1308 7352 1360 7404
rect 2780 7352 2832 7404
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 9680 7352 9732 7404
rect 3516 7284 3568 7336
rect 3608 7191 3660 7200
rect 3608 7157 3617 7191
rect 3617 7157 3651 7191
rect 3651 7157 3660 7191
rect 3608 7148 3660 7157
rect 10048 7191 10100 7200
rect 10048 7157 10057 7191
rect 10057 7157 10091 7191
rect 10091 7157 10100 7191
rect 10048 7148 10100 7157
rect 2582 7046 2634 7098
rect 2646 7046 2698 7098
rect 2710 7046 2762 7098
rect 2774 7046 2826 7098
rect 2838 7046 2890 7098
rect 5845 7046 5897 7098
rect 5909 7046 5961 7098
rect 5973 7046 6025 7098
rect 6037 7046 6089 7098
rect 6101 7046 6153 7098
rect 9109 7046 9161 7098
rect 9173 7046 9225 7098
rect 9237 7046 9289 7098
rect 9301 7046 9353 7098
rect 9365 7046 9417 7098
rect 3608 6944 3660 6996
rect 9772 6944 9824 6996
rect 3056 6808 3108 6860
rect 2872 6740 2924 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 1860 6715 1912 6724
rect 1860 6681 1869 6715
rect 1869 6681 1903 6715
rect 1903 6681 1912 6715
rect 1860 6672 1912 6681
rect 6460 6672 6512 6724
rect 2872 6604 2924 6656
rect 3056 6604 3108 6656
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 10048 6647 10100 6656
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 4213 6502 4265 6554
rect 4277 6502 4329 6554
rect 4341 6502 4393 6554
rect 4405 6502 4457 6554
rect 4469 6502 4521 6554
rect 7477 6502 7529 6554
rect 7541 6502 7593 6554
rect 7605 6502 7657 6554
rect 7669 6502 7721 6554
rect 7733 6502 7785 6554
rect 4068 6400 4120 6452
rect 2044 6264 2096 6316
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 3884 6196 3936 6248
rect 9864 6128 9916 6180
rect 4804 6060 4856 6112
rect 2582 5958 2634 6010
rect 2646 5958 2698 6010
rect 2710 5958 2762 6010
rect 2774 5958 2826 6010
rect 2838 5958 2890 6010
rect 5845 5958 5897 6010
rect 5909 5958 5961 6010
rect 5973 5958 6025 6010
rect 6037 5958 6089 6010
rect 6101 5958 6153 6010
rect 9109 5958 9161 6010
rect 9173 5958 9225 6010
rect 9237 5958 9289 6010
rect 9301 5958 9353 6010
rect 9365 5958 9417 6010
rect 2964 5856 3016 5908
rect 3332 5856 3384 5908
rect 6828 5788 6880 5840
rect 9680 5788 9732 5840
rect 2044 5652 2096 5704
rect 3056 5720 3108 5772
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 9680 5652 9732 5704
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 4213 5414 4265 5466
rect 4277 5414 4329 5466
rect 4341 5414 4393 5466
rect 4405 5414 4457 5466
rect 4469 5414 4521 5466
rect 7477 5414 7529 5466
rect 7541 5414 7593 5466
rect 7605 5414 7657 5466
rect 7669 5414 7721 5466
rect 7733 5414 7785 5466
rect 3516 5312 3568 5364
rect 1216 5244 1268 5296
rect 3240 5176 3292 5228
rect 3516 5176 3568 5228
rect 3332 5108 3384 5160
rect 6368 4972 6420 5024
rect 10048 5015 10100 5024
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 2582 4870 2634 4922
rect 2646 4870 2698 4922
rect 2710 4870 2762 4922
rect 2774 4870 2826 4922
rect 2838 4870 2890 4922
rect 5845 4870 5897 4922
rect 5909 4870 5961 4922
rect 5973 4870 6025 4922
rect 6037 4870 6089 4922
rect 6101 4870 6153 4922
rect 9109 4870 9161 4922
rect 9173 4870 9225 4922
rect 9237 4870 9289 4922
rect 9301 4870 9353 4922
rect 9365 4870 9417 4922
rect 3148 4768 3200 4820
rect 6276 4700 6328 4752
rect 1584 4564 1636 4616
rect 1676 4496 1728 4548
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 9772 4564 9824 4616
rect 9680 4496 9732 4548
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 10048 4471 10100 4480
rect 10048 4437 10057 4471
rect 10057 4437 10091 4471
rect 10091 4437 10100 4471
rect 10048 4428 10100 4437
rect 4213 4326 4265 4378
rect 4277 4326 4329 4378
rect 4341 4326 4393 4378
rect 4405 4326 4457 4378
rect 4469 4326 4521 4378
rect 7477 4326 7529 4378
rect 7541 4326 7593 4378
rect 7605 4326 7657 4378
rect 7669 4326 7721 4378
rect 7733 4326 7785 4378
rect 3240 4224 3292 4276
rect 9772 4224 9824 4276
rect 1216 4088 1268 4140
rect 2228 4088 2280 4140
rect 2504 4088 2556 4140
rect 3516 4131 3568 4140
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 3608 4088 3660 4140
rect 5540 4020 5592 4072
rect 9864 3952 9916 4004
rect 3056 3884 3108 3936
rect 2582 3782 2634 3834
rect 2646 3782 2698 3834
rect 2710 3782 2762 3834
rect 2774 3782 2826 3834
rect 2838 3782 2890 3834
rect 5845 3782 5897 3834
rect 5909 3782 5961 3834
rect 5973 3782 6025 3834
rect 6037 3782 6089 3834
rect 6101 3782 6153 3834
rect 9109 3782 9161 3834
rect 9173 3782 9225 3834
rect 9237 3782 9289 3834
rect 9301 3782 9353 3834
rect 9365 3782 9417 3834
rect 2320 3680 2372 3732
rect 8116 3612 8168 3664
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2412 3476 2464 3528
rect 3516 3476 3568 3528
rect 3792 3408 3844 3460
rect 10048 3383 10100 3392
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 4213 3238 4265 3290
rect 4277 3238 4329 3290
rect 4341 3238 4393 3290
rect 4405 3238 4457 3290
rect 4469 3238 4521 3290
rect 7477 3238 7529 3290
rect 7541 3238 7593 3290
rect 7605 3238 7657 3290
rect 7669 3238 7721 3290
rect 7733 3238 7785 3290
rect 2228 3136 2280 3188
rect 2136 3000 2188 3052
rect 2872 3043 2924 3052
rect 2872 3009 2881 3043
rect 2881 3009 2915 3043
rect 2915 3009 2924 3043
rect 2872 3000 2924 3009
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 3608 3000 3660 3052
rect 6368 3000 6420 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 2044 2864 2096 2916
rect 3332 2907 3384 2916
rect 3332 2873 3341 2907
rect 3341 2873 3375 2907
rect 3375 2873 3384 2907
rect 3332 2864 3384 2873
rect 9496 2796 9548 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 2582 2694 2634 2746
rect 2646 2694 2698 2746
rect 2710 2694 2762 2746
rect 2774 2694 2826 2746
rect 2838 2694 2890 2746
rect 5845 2694 5897 2746
rect 5909 2694 5961 2746
rect 5973 2694 6025 2746
rect 6037 2694 6089 2746
rect 6101 2694 6153 2746
rect 9109 2694 9161 2746
rect 9173 2694 9225 2746
rect 9237 2694 9289 2746
rect 9301 2694 9353 2746
rect 9365 2694 9417 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 1676 2592 1728 2644
rect 2504 2592 2556 2644
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 3884 2592 3936 2644
rect 1308 2388 1360 2440
rect 2780 2388 2832 2440
rect 2872 2431 2924 2440
rect 2872 2397 2881 2431
rect 2881 2397 2915 2431
rect 2915 2397 2924 2431
rect 3976 2431 4028 2440
rect 2872 2388 2924 2397
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 9036 2388 9088 2440
rect 9772 2388 9824 2440
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 10048 2295 10100 2304
rect 10048 2261 10057 2295
rect 10057 2261 10091 2295
rect 10091 2261 10100 2295
rect 10048 2252 10100 2261
rect 4213 2150 4265 2202
rect 4277 2150 4329 2202
rect 4341 2150 4393 2202
rect 4405 2150 4457 2202
rect 4469 2150 4521 2202
rect 7477 2150 7529 2202
rect 7541 2150 7593 2202
rect 7605 2150 7657 2202
rect 7669 2150 7721 2202
rect 7733 2150 7785 2202
rect 2780 484 2832 536
rect 4620 484 4672 536
<< metal2 >>
rect 2962 79656 3018 79665
rect 2962 79591 3018 79600
rect 2582 77820 2890 77840
rect 2582 77818 2588 77820
rect 2644 77818 2668 77820
rect 2724 77818 2748 77820
rect 2804 77818 2828 77820
rect 2884 77818 2890 77820
rect 2644 77766 2646 77818
rect 2826 77766 2828 77818
rect 2582 77764 2588 77766
rect 2644 77764 2668 77766
rect 2724 77764 2748 77766
rect 2804 77764 2828 77766
rect 2884 77764 2890 77766
rect 2582 77744 2890 77764
rect 2504 77512 2556 77518
rect 2504 77454 2556 77460
rect 1124 77444 1176 77450
rect 1124 77386 1176 77392
rect 388 75472 440 75478
rect 388 75414 440 75420
rect 204 50788 256 50794
rect 204 50730 256 50736
rect 112 50516 164 50522
rect 112 50458 164 50464
rect 124 44062 152 50458
rect 216 48210 244 50730
rect 296 49768 348 49774
rect 296 49710 348 49716
rect 204 48204 256 48210
rect 204 48146 256 48152
rect 112 44056 164 44062
rect 112 43998 164 44004
rect 216 36582 244 48146
rect 204 36576 256 36582
rect 204 36518 256 36524
rect 308 30734 336 49710
rect 400 48346 428 75414
rect 940 70372 992 70378
rect 940 70314 992 70320
rect 480 65476 532 65482
rect 480 65418 532 65424
rect 388 48340 440 48346
rect 388 48282 440 48288
rect 388 48068 440 48074
rect 388 48010 440 48016
rect 296 30728 348 30734
rect 296 30670 348 30676
rect 400 28762 428 48010
rect 492 46034 520 65418
rect 952 62830 980 70314
rect 1032 65544 1084 65550
rect 1032 65486 1084 65492
rect 940 62824 992 62830
rect 940 62766 992 62772
rect 664 62484 716 62490
rect 664 62426 716 62432
rect 572 52080 624 52086
rect 572 52022 624 52028
rect 480 46028 532 46034
rect 480 45970 532 45976
rect 388 28756 440 28762
rect 388 28698 440 28704
rect 584 24750 612 52022
rect 676 49434 704 62426
rect 940 59696 992 59702
rect 940 59638 992 59644
rect 848 59424 900 59430
rect 848 59366 900 59372
rect 756 59016 808 59022
rect 756 58958 808 58964
rect 664 49428 716 49434
rect 664 49370 716 49376
rect 664 48816 716 48822
rect 664 48758 716 48764
rect 676 44198 704 48758
rect 664 44192 716 44198
rect 664 44134 716 44140
rect 664 44056 716 44062
rect 664 43998 716 44004
rect 676 27062 704 43998
rect 768 40186 796 58958
rect 860 58857 888 59366
rect 846 58848 902 58857
rect 846 58783 902 58792
rect 848 58540 900 58546
rect 848 58482 900 58488
rect 756 40180 808 40186
rect 756 40122 808 40128
rect 860 39030 888 58482
rect 952 43450 980 59638
rect 1044 44946 1072 65486
rect 1136 57798 1164 77386
rect 2516 77081 2544 77454
rect 2976 77450 3004 79591
rect 3882 79248 3938 79257
rect 3882 79183 3938 79192
rect 3054 78840 3110 78849
rect 3054 78775 3110 78784
rect 3068 77586 3096 78775
rect 3330 78432 3386 78441
rect 3330 78367 3386 78376
rect 3240 77648 3292 77654
rect 3240 77590 3292 77596
rect 3056 77580 3108 77586
rect 3056 77522 3108 77528
rect 2964 77444 3016 77450
rect 2964 77386 3016 77392
rect 3056 77376 3108 77382
rect 3056 77318 3108 77324
rect 2502 77072 2558 77081
rect 1400 77036 1452 77042
rect 1400 76978 1452 76984
rect 2044 77036 2096 77042
rect 2502 77007 2558 77016
rect 2780 77036 2832 77042
rect 2044 76978 2096 76984
rect 2780 76978 2832 76984
rect 1216 76560 1268 76566
rect 1216 76502 1268 76508
rect 1124 57792 1176 57798
rect 1124 57734 1176 57740
rect 1124 57520 1176 57526
rect 1122 57488 1124 57497
rect 1176 57488 1178 57497
rect 1122 57423 1178 57432
rect 1228 55876 1256 76502
rect 1412 75449 1440 76978
rect 1584 76832 1636 76838
rect 1584 76774 1636 76780
rect 1398 75440 1454 75449
rect 1398 75375 1454 75384
rect 1308 75336 1360 75342
rect 1308 75278 1360 75284
rect 1320 74089 1348 75278
rect 1400 74860 1452 74866
rect 1400 74802 1452 74808
rect 1306 74080 1362 74089
rect 1306 74015 1362 74024
rect 1412 73681 1440 74802
rect 1596 74254 1624 76774
rect 1860 76628 1912 76634
rect 1860 76570 1912 76576
rect 1676 76424 1728 76430
rect 1676 76366 1728 76372
rect 1688 75954 1716 76366
rect 1872 76022 1900 76570
rect 2056 76265 2084 76978
rect 2792 76945 2820 76978
rect 2778 76936 2834 76945
rect 2778 76871 2834 76880
rect 2228 76832 2280 76838
rect 2228 76774 2280 76780
rect 2136 76424 2188 76430
rect 2136 76366 2188 76372
rect 2042 76256 2098 76265
rect 2042 76191 2098 76200
rect 1860 76016 1912 76022
rect 1860 75958 1912 75964
rect 2148 75954 2176 76366
rect 1676 75948 1728 75954
rect 1676 75890 1728 75896
rect 2136 75948 2188 75954
rect 2136 75890 2188 75896
rect 1768 75744 1820 75750
rect 1768 75686 1820 75692
rect 1584 74248 1636 74254
rect 1584 74190 1636 74196
rect 1492 74180 1544 74186
rect 1492 74122 1544 74128
rect 1504 73778 1532 74122
rect 1492 73772 1544 73778
rect 1492 73714 1544 73720
rect 1398 73672 1454 73681
rect 1398 73607 1454 73616
rect 1400 73160 1452 73166
rect 1400 73102 1452 73108
rect 1308 72684 1360 72690
rect 1308 72626 1360 72632
rect 1320 71913 1348 72626
rect 1412 72457 1440 73102
rect 1398 72448 1454 72457
rect 1398 72383 1454 72392
rect 1400 72276 1452 72282
rect 1400 72218 1452 72224
rect 1412 72078 1440 72218
rect 1400 72072 1452 72078
rect 1400 72014 1452 72020
rect 1306 71904 1362 71913
rect 1306 71839 1362 71848
rect 1412 71618 1440 72014
rect 1504 71942 1532 73714
rect 1676 73024 1728 73030
rect 1676 72966 1728 72972
rect 1492 71936 1544 71942
rect 1492 71878 1544 71884
rect 1412 71590 1624 71618
rect 1400 71528 1452 71534
rect 1306 71496 1362 71505
rect 1400 71470 1452 71476
rect 1306 71431 1362 71440
rect 1320 71058 1348 71431
rect 1412 71097 1440 71470
rect 1398 71088 1454 71097
rect 1308 71052 1360 71058
rect 1398 71023 1454 71032
rect 1308 70994 1360 71000
rect 1596 70310 1624 71590
rect 1584 70304 1636 70310
rect 1306 70272 1362 70281
rect 1584 70246 1636 70252
rect 1306 70207 1362 70216
rect 1320 69902 1348 70207
rect 1308 69896 1360 69902
rect 1308 69838 1360 69844
rect 1596 69737 1624 70246
rect 1582 69728 1638 69737
rect 1582 69663 1638 69672
rect 1584 69556 1636 69562
rect 1584 69498 1636 69504
rect 1596 69426 1624 69498
rect 1584 69420 1636 69426
rect 1584 69362 1636 69368
rect 1688 69306 1716 72966
rect 1780 72185 1808 75686
rect 1860 75200 1912 75206
rect 1860 75142 1912 75148
rect 1766 72176 1822 72185
rect 1766 72111 1822 72120
rect 1768 72072 1820 72078
rect 1768 72014 1820 72020
rect 1780 71942 1808 72014
rect 1768 71936 1820 71942
rect 1768 71878 1820 71884
rect 1768 71528 1820 71534
rect 1768 71470 1820 71476
rect 1780 70378 1808 71470
rect 1768 70372 1820 70378
rect 1768 70314 1820 70320
rect 1768 69488 1820 69494
rect 1766 69456 1768 69465
rect 1820 69456 1822 69465
rect 1766 69391 1822 69400
rect 1400 69284 1452 69290
rect 1400 69226 1452 69232
rect 1596 69278 1716 69306
rect 1768 69352 1820 69358
rect 1768 69294 1820 69300
rect 1308 68808 1360 68814
rect 1308 68750 1360 68756
rect 1320 67697 1348 68750
rect 1412 67862 1440 69226
rect 1492 69216 1544 69222
rect 1492 69158 1544 69164
rect 1504 69057 1532 69158
rect 1490 69048 1546 69057
rect 1490 68983 1546 68992
rect 1492 68264 1544 68270
rect 1492 68206 1544 68212
rect 1400 67856 1452 67862
rect 1400 67798 1452 67804
rect 1400 67720 1452 67726
rect 1306 67688 1362 67697
rect 1400 67662 1452 67668
rect 1306 67623 1362 67632
rect 1412 67289 1440 67662
rect 1398 67280 1454 67289
rect 1504 67250 1532 68206
rect 1398 67215 1454 67224
rect 1492 67244 1544 67250
rect 1492 67186 1544 67192
rect 1504 66586 1532 67186
rect 1412 66558 1532 66586
rect 1412 66178 1440 66558
rect 1492 66496 1544 66502
rect 1492 66438 1544 66444
rect 1320 66150 1440 66178
rect 1320 65770 1348 66150
rect 1400 66088 1452 66094
rect 1400 66030 1452 66036
rect 1412 65929 1440 66030
rect 1398 65920 1454 65929
rect 1398 65855 1454 65864
rect 1320 65742 1440 65770
rect 1412 65006 1440 65742
rect 1504 65521 1532 66438
rect 1490 65512 1546 65521
rect 1490 65447 1546 65456
rect 1492 65408 1544 65414
rect 1492 65350 1544 65356
rect 1400 65000 1452 65006
rect 1400 64942 1452 64948
rect 1400 64320 1452 64326
rect 1504 64297 1532 65350
rect 1400 64262 1452 64268
rect 1490 64288 1546 64297
rect 1412 62529 1440 64262
rect 1490 64223 1546 64232
rect 1596 63918 1624 69278
rect 1676 68332 1728 68338
rect 1676 68274 1728 68280
rect 1688 67182 1716 68274
rect 1676 67176 1728 67182
rect 1676 67118 1728 67124
rect 1688 65074 1716 67118
rect 1676 65068 1728 65074
rect 1676 65010 1728 65016
rect 1688 64598 1716 65010
rect 1676 64592 1728 64598
rect 1676 64534 1728 64540
rect 1584 63912 1636 63918
rect 1584 63854 1636 63860
rect 1688 63442 1716 64534
rect 1676 63436 1728 63442
rect 1676 63378 1728 63384
rect 1676 63300 1728 63306
rect 1676 63242 1728 63248
rect 1688 63034 1716 63242
rect 1676 63028 1728 63034
rect 1676 62970 1728 62976
rect 1584 62892 1636 62898
rect 1584 62834 1636 62840
rect 1492 62688 1544 62694
rect 1492 62630 1544 62636
rect 1398 62520 1454 62529
rect 1398 62455 1454 62464
rect 1400 62416 1452 62422
rect 1400 62358 1452 62364
rect 1412 60858 1440 62358
rect 1504 61713 1532 62630
rect 1490 61704 1546 61713
rect 1490 61639 1546 61648
rect 1596 60874 1624 62834
rect 1780 62422 1808 69294
rect 1872 68474 1900 75142
rect 1952 74656 2004 74662
rect 1952 74598 2004 74604
rect 1860 68468 1912 68474
rect 1860 68410 1912 68416
rect 1964 68406 1992 74598
rect 2136 74112 2188 74118
rect 2136 74054 2188 74060
rect 2148 73778 2176 74054
rect 2136 73772 2188 73778
rect 2136 73714 2188 73720
rect 2044 73024 2096 73030
rect 2044 72966 2096 72972
rect 1952 68400 2004 68406
rect 1952 68342 2004 68348
rect 1860 67720 1912 67726
rect 2056 67674 2084 72966
rect 2148 72282 2176 73714
rect 2240 73658 2268 76774
rect 2582 76732 2890 76752
rect 2582 76730 2588 76732
rect 2644 76730 2668 76732
rect 2724 76730 2748 76732
rect 2804 76730 2828 76732
rect 2884 76730 2890 76732
rect 2644 76678 2646 76730
rect 2826 76678 2828 76730
rect 2582 76676 2588 76678
rect 2644 76676 2668 76678
rect 2724 76676 2748 76678
rect 2804 76676 2828 76678
rect 2884 76676 2890 76678
rect 2582 76656 2890 76676
rect 2780 76560 2832 76566
rect 2780 76502 2832 76508
rect 2792 76430 2820 76502
rect 2780 76424 2832 76430
rect 2780 76366 2832 76372
rect 2964 76424 3016 76430
rect 2964 76366 3016 76372
rect 2976 75857 3004 76366
rect 2962 75848 3018 75857
rect 2962 75783 3018 75792
rect 2582 75644 2890 75664
rect 2582 75642 2588 75644
rect 2644 75642 2668 75644
rect 2724 75642 2748 75644
rect 2804 75642 2828 75644
rect 2884 75642 2890 75644
rect 2644 75590 2646 75642
rect 2826 75590 2828 75642
rect 2582 75588 2588 75590
rect 2644 75588 2668 75590
rect 2724 75588 2748 75590
rect 2804 75588 2828 75590
rect 2884 75588 2890 75590
rect 2582 75568 2890 75588
rect 2596 75336 2648 75342
rect 2596 75278 2648 75284
rect 2964 75336 3016 75342
rect 2964 75278 3016 75284
rect 2608 74866 2636 75278
rect 2872 74996 2924 75002
rect 2872 74938 2924 74944
rect 2884 74866 2912 74938
rect 2976 74866 3004 75278
rect 3068 75206 3096 77318
rect 3148 76288 3200 76294
rect 3148 76230 3200 76236
rect 3056 75200 3108 75206
rect 3056 75142 3108 75148
rect 2596 74860 2648 74866
rect 2596 74802 2648 74808
rect 2872 74860 2924 74866
rect 2872 74802 2924 74808
rect 2964 74860 3016 74866
rect 2964 74802 3016 74808
rect 2608 74746 2636 74802
rect 2516 74718 2636 74746
rect 2516 74254 2544 74718
rect 2582 74556 2890 74576
rect 2582 74554 2588 74556
rect 2644 74554 2668 74556
rect 2724 74554 2748 74556
rect 2804 74554 2828 74556
rect 2884 74554 2890 74556
rect 2644 74502 2646 74554
rect 2826 74502 2828 74554
rect 2582 74500 2588 74502
rect 2644 74500 2668 74502
rect 2724 74500 2748 74502
rect 2804 74500 2828 74502
rect 2884 74500 2890 74502
rect 2582 74480 2890 74500
rect 2504 74248 2556 74254
rect 2504 74190 2556 74196
rect 2780 74248 2832 74254
rect 2780 74190 2832 74196
rect 2792 73930 2820 74190
rect 2792 73902 3096 73930
rect 2964 73772 3016 73778
rect 2964 73714 3016 73720
rect 2240 73630 2452 73658
rect 2320 73568 2372 73574
rect 2320 73510 2372 73516
rect 2228 73160 2280 73166
rect 2228 73102 2280 73108
rect 2240 72865 2268 73102
rect 2226 72856 2282 72865
rect 2226 72791 2282 72800
rect 2228 72480 2280 72486
rect 2228 72422 2280 72428
rect 2136 72276 2188 72282
rect 2136 72218 2188 72224
rect 2134 72176 2190 72185
rect 2134 72111 2190 72120
rect 2148 69494 2176 72111
rect 2136 69488 2188 69494
rect 2136 69430 2188 69436
rect 2136 68672 2188 68678
rect 2136 68614 2188 68620
rect 1860 67662 1912 67668
rect 1768 62416 1820 62422
rect 1768 62358 1820 62364
rect 1768 62280 1820 62286
rect 1768 62222 1820 62228
rect 1780 61810 1808 62222
rect 1768 61804 1820 61810
rect 1768 61746 1820 61752
rect 1780 61690 1808 61746
rect 1688 61662 1808 61690
rect 1688 61198 1716 61662
rect 1768 61396 1820 61402
rect 1768 61338 1820 61344
rect 1676 61192 1728 61198
rect 1676 61134 1728 61140
rect 1400 60852 1452 60858
rect 1400 60794 1452 60800
rect 1504 60846 1624 60874
rect 1504 60734 1532 60846
rect 1320 60722 1532 60734
rect 1584 60784 1636 60790
rect 1584 60726 1636 60732
rect 1308 60716 1532 60722
rect 1360 60706 1532 60716
rect 1308 60658 1360 60664
rect 1492 60512 1544 60518
rect 1492 60454 1544 60460
rect 1308 59968 1360 59974
rect 1504 59945 1532 60454
rect 1308 59910 1360 59916
rect 1490 59936 1546 59945
rect 1320 59129 1348 59910
rect 1490 59871 1546 59880
rect 1492 59628 1544 59634
rect 1492 59570 1544 59576
rect 1400 59560 1452 59566
rect 1398 59528 1400 59537
rect 1452 59528 1454 59537
rect 1398 59463 1454 59472
rect 1306 59120 1362 59129
rect 1306 59055 1362 59064
rect 1504 58970 1532 59570
rect 1320 58942 1532 58970
rect 1320 57905 1348 58942
rect 1492 58880 1544 58886
rect 1492 58822 1544 58828
rect 1400 58336 1452 58342
rect 1400 58278 1452 58284
rect 1306 57896 1362 57905
rect 1306 57831 1362 57840
rect 1308 57792 1360 57798
rect 1308 57734 1360 57740
rect 1320 56386 1348 57734
rect 1412 57361 1440 58278
rect 1504 58177 1532 58822
rect 1490 58168 1546 58177
rect 1490 58103 1546 58112
rect 1492 57996 1544 58002
rect 1492 57938 1544 57944
rect 1504 57458 1532 57938
rect 1492 57452 1544 57458
rect 1492 57394 1544 57400
rect 1398 57352 1454 57361
rect 1398 57287 1454 57296
rect 1398 56944 1454 56953
rect 1398 56879 1454 56888
rect 1412 56506 1440 56879
rect 1492 56704 1544 56710
rect 1492 56646 1544 56652
rect 1504 56545 1532 56646
rect 1490 56536 1546 56545
rect 1400 56500 1452 56506
rect 1490 56471 1546 56480
rect 1400 56442 1452 56448
rect 1320 56358 1440 56386
rect 1136 55848 1256 55876
rect 1032 44940 1084 44946
rect 1032 44882 1084 44888
rect 1136 44538 1164 55848
rect 1412 52986 1440 56358
rect 1492 55616 1544 55622
rect 1492 55558 1544 55564
rect 1504 54777 1532 55558
rect 1490 54768 1546 54777
rect 1490 54703 1546 54712
rect 1492 54528 1544 54534
rect 1492 54470 1544 54476
rect 1504 53961 1532 54470
rect 1490 53952 1546 53961
rect 1490 53887 1546 53896
rect 1492 53576 1544 53582
rect 1492 53518 1544 53524
rect 1504 53242 1532 53518
rect 1492 53236 1544 53242
rect 1492 53178 1544 53184
rect 1320 52958 1440 52986
rect 1216 52488 1268 52494
rect 1216 52430 1268 52436
rect 1228 50402 1256 52430
rect 1320 52068 1348 52958
rect 1400 52896 1452 52902
rect 1400 52838 1452 52844
rect 1412 52193 1440 52838
rect 1492 52352 1544 52358
rect 1492 52294 1544 52300
rect 1398 52184 1454 52193
rect 1398 52119 1454 52128
rect 1320 52040 1440 52068
rect 1308 51808 1360 51814
rect 1308 51750 1360 51756
rect 1320 51097 1348 51750
rect 1412 51626 1440 52040
rect 1504 51785 1532 52294
rect 1490 51776 1546 51785
rect 1490 51711 1546 51720
rect 1412 51598 1532 51626
rect 1400 51264 1452 51270
rect 1400 51206 1452 51212
rect 1306 51088 1362 51097
rect 1306 51023 1362 51032
rect 1412 50912 1440 51206
rect 1320 50884 1440 50912
rect 1320 50561 1348 50884
rect 1504 50810 1532 51598
rect 1412 50782 1532 50810
rect 1306 50552 1362 50561
rect 1306 50487 1362 50496
rect 1228 50374 1348 50402
rect 1216 50244 1268 50250
rect 1216 50186 1268 50192
rect 1124 44532 1176 44538
rect 1124 44474 1176 44480
rect 1124 44192 1176 44198
rect 1124 44134 1176 44140
rect 940 43444 992 43450
rect 940 43386 992 43392
rect 1032 41540 1084 41546
rect 1032 41482 1084 41488
rect 848 39024 900 39030
rect 848 38966 900 38972
rect 940 36576 992 36582
rect 940 36518 992 36524
rect 952 31414 980 36518
rect 940 31408 992 31414
rect 940 31350 992 31356
rect 664 27056 716 27062
rect 664 26998 716 27004
rect 572 24744 624 24750
rect 572 24686 624 24692
rect 1044 23798 1072 41482
rect 1136 25498 1164 44134
rect 1228 32910 1256 50186
rect 1320 43636 1348 50374
rect 1412 49230 1440 50782
rect 1492 50720 1544 50726
rect 1492 50662 1544 50668
rect 1504 50017 1532 50662
rect 1596 50318 1624 60726
rect 1688 60246 1716 61134
rect 1676 60240 1728 60246
rect 1676 60182 1728 60188
rect 1676 59764 1728 59770
rect 1676 59706 1728 59712
rect 1688 57594 1716 59706
rect 1676 57588 1728 57594
rect 1676 57530 1728 57536
rect 1676 57248 1728 57254
rect 1676 57190 1728 57196
rect 1688 56846 1716 57190
rect 1676 56840 1728 56846
rect 1676 56782 1728 56788
rect 1676 56500 1728 56506
rect 1676 56442 1728 56448
rect 1688 55214 1716 56442
rect 1676 55208 1728 55214
rect 1676 55150 1728 55156
rect 1676 55072 1728 55078
rect 1676 55014 1728 55020
rect 1688 54126 1716 55014
rect 1676 54120 1728 54126
rect 1676 54062 1728 54068
rect 1688 53242 1716 54062
rect 1780 53718 1808 61338
rect 1872 60858 1900 67662
rect 1964 67646 2084 67674
rect 1964 65142 1992 67646
rect 2148 66586 2176 68614
rect 2056 66558 2176 66586
rect 1952 65136 2004 65142
rect 1952 65078 2004 65084
rect 1952 65000 2004 65006
rect 1952 64942 2004 64948
rect 1964 63986 1992 64942
rect 1952 63980 2004 63986
rect 1952 63922 2004 63928
rect 1964 63374 1992 63922
rect 1952 63368 2004 63374
rect 1952 63310 2004 63316
rect 1952 62144 2004 62150
rect 1952 62086 2004 62092
rect 1964 61606 1992 62086
rect 2056 61985 2084 66558
rect 2136 66496 2188 66502
rect 2136 66438 2188 66444
rect 2042 61976 2098 61985
rect 2042 61911 2098 61920
rect 2044 61804 2096 61810
rect 2044 61746 2096 61752
rect 1952 61600 2004 61606
rect 1952 61542 2004 61548
rect 1964 61266 1992 61542
rect 1952 61260 2004 61266
rect 1952 61202 2004 61208
rect 1860 60852 1912 60858
rect 1860 60794 1912 60800
rect 1860 60716 1912 60722
rect 1860 60658 1912 60664
rect 1872 60314 1900 60658
rect 1860 60308 1912 60314
rect 1860 60250 1912 60256
rect 1964 60194 1992 61202
rect 1872 60166 1992 60194
rect 1872 59090 1900 60166
rect 1952 60104 2004 60110
rect 1952 60046 2004 60052
rect 1860 59084 1912 59090
rect 1860 59026 1912 59032
rect 1872 58070 1900 59026
rect 1860 58064 1912 58070
rect 1860 58006 1912 58012
rect 1964 57934 1992 60046
rect 1952 57928 2004 57934
rect 1858 57896 1914 57905
rect 1952 57870 2004 57876
rect 1858 57831 1914 57840
rect 1872 56438 1900 57831
rect 1964 57458 1992 57870
rect 1952 57452 2004 57458
rect 1952 57394 2004 57400
rect 1860 56432 1912 56438
rect 1860 56374 1912 56380
rect 1860 56228 1912 56234
rect 1860 56170 1912 56176
rect 1872 55282 1900 56170
rect 2056 55706 2084 61746
rect 2148 61402 2176 66438
rect 2240 66178 2268 72422
rect 2332 67250 2360 73510
rect 2424 69834 2452 73630
rect 2582 73468 2890 73488
rect 2582 73466 2588 73468
rect 2644 73466 2668 73468
rect 2724 73466 2748 73468
rect 2804 73466 2828 73468
rect 2884 73466 2890 73468
rect 2644 73414 2646 73466
rect 2826 73414 2828 73466
rect 2582 73412 2588 73414
rect 2644 73412 2668 73414
rect 2724 73412 2748 73414
rect 2804 73412 2828 73414
rect 2884 73412 2890 73414
rect 2582 73392 2890 73412
rect 2976 73273 3004 73714
rect 2962 73264 3018 73273
rect 2962 73199 3018 73208
rect 2582 72380 2890 72400
rect 2582 72378 2588 72380
rect 2644 72378 2668 72380
rect 2724 72378 2748 72380
rect 2804 72378 2828 72380
rect 2884 72378 2890 72380
rect 2644 72326 2646 72378
rect 2826 72326 2828 72378
rect 2582 72324 2588 72326
rect 2644 72324 2668 72326
rect 2724 72324 2748 72326
rect 2804 72324 2828 72326
rect 2884 72324 2890 72326
rect 2582 72304 2890 72324
rect 2582 71292 2890 71312
rect 2582 71290 2588 71292
rect 2644 71290 2668 71292
rect 2724 71290 2748 71292
rect 2804 71290 2828 71292
rect 2884 71290 2890 71292
rect 2644 71238 2646 71290
rect 2826 71238 2828 71290
rect 2582 71236 2588 71238
rect 2644 71236 2668 71238
rect 2724 71236 2748 71238
rect 2804 71236 2828 71238
rect 2884 71236 2890 71238
rect 2582 71216 2890 71236
rect 2504 70984 2556 70990
rect 2504 70926 2556 70932
rect 2780 70984 2832 70990
rect 2780 70926 2832 70932
rect 2412 69828 2464 69834
rect 2412 69770 2464 69776
rect 2410 69728 2466 69737
rect 2410 69663 2466 69672
rect 2424 69426 2452 69663
rect 2412 69420 2464 69426
rect 2412 69362 2464 69368
rect 2424 68338 2452 69362
rect 2412 68332 2464 68338
rect 2412 68274 2464 68280
rect 2320 67244 2372 67250
rect 2320 67186 2372 67192
rect 2320 66632 2372 66638
rect 2320 66574 2372 66580
rect 2332 66337 2360 66574
rect 2318 66328 2374 66337
rect 2318 66263 2374 66272
rect 2240 66150 2452 66178
rect 2320 65408 2372 65414
rect 2320 65350 2372 65356
rect 2332 64841 2360 65350
rect 2318 64832 2374 64841
rect 2318 64767 2374 64776
rect 2424 64682 2452 66150
rect 2332 64654 2452 64682
rect 2332 63238 2360 64654
rect 2412 64524 2464 64530
rect 2412 64466 2464 64472
rect 2424 63986 2452 64466
rect 2412 63980 2464 63986
rect 2412 63922 2464 63928
rect 2412 63368 2464 63374
rect 2412 63310 2464 63316
rect 2320 63232 2372 63238
rect 2320 63174 2372 63180
rect 2320 62960 2372 62966
rect 2424 62948 2452 63310
rect 2372 62920 2452 62948
rect 2320 62902 2372 62908
rect 2320 62824 2372 62830
rect 2320 62766 2372 62772
rect 2228 62688 2280 62694
rect 2228 62630 2280 62636
rect 2240 62121 2268 62630
rect 2226 62112 2282 62121
rect 2226 62047 2282 62056
rect 2226 61976 2282 61985
rect 2226 61911 2282 61920
rect 2136 61396 2188 61402
rect 2136 61338 2188 61344
rect 2240 61282 2268 61911
rect 2148 61254 2268 61282
rect 2148 57798 2176 61254
rect 2228 61192 2280 61198
rect 2228 61134 2280 61140
rect 2136 57792 2188 57798
rect 2136 57734 2188 57740
rect 2136 57588 2188 57594
rect 2136 57530 2188 57536
rect 1964 55678 2084 55706
rect 1860 55276 1912 55282
rect 1860 55218 1912 55224
rect 1768 53712 1820 53718
rect 1768 53654 1820 53660
rect 1872 53582 1900 55218
rect 1860 53576 1912 53582
rect 1860 53518 1912 53524
rect 1768 53440 1820 53446
rect 1768 53382 1820 53388
rect 1676 53236 1728 53242
rect 1676 53178 1728 53184
rect 1676 51808 1728 51814
rect 1676 51750 1728 51756
rect 1688 51406 1716 51750
rect 1676 51400 1728 51406
rect 1676 51342 1728 51348
rect 1676 51264 1728 51270
rect 1676 51206 1728 51212
rect 1688 50522 1716 51206
rect 1676 50516 1728 50522
rect 1676 50458 1728 50464
rect 1676 50380 1728 50386
rect 1676 50322 1728 50328
rect 1584 50312 1636 50318
rect 1584 50254 1636 50260
rect 1584 50176 1636 50182
rect 1584 50118 1636 50124
rect 1490 50008 1546 50017
rect 1490 49943 1546 49952
rect 1596 49586 1624 50118
rect 1688 49774 1716 50322
rect 1780 49978 1808 53382
rect 1872 50318 1900 53518
rect 1964 51048 1992 55678
rect 2148 53446 2176 57530
rect 2240 54641 2268 61134
rect 2332 60636 2360 62766
rect 2424 62286 2452 62920
rect 2412 62280 2464 62286
rect 2412 62222 2464 62228
rect 2424 60858 2452 62222
rect 2412 60852 2464 60858
rect 2412 60794 2464 60800
rect 2332 60608 2452 60636
rect 2320 60512 2372 60518
rect 2320 60454 2372 60460
rect 2332 57458 2360 60454
rect 2424 57594 2452 60608
rect 2516 59786 2544 70926
rect 2792 70689 2820 70926
rect 2778 70680 2834 70689
rect 2688 70644 2740 70650
rect 2778 70615 2834 70624
rect 2872 70644 2924 70650
rect 2688 70586 2740 70592
rect 2872 70586 2924 70592
rect 2700 70394 2728 70586
rect 2884 70530 2912 70586
rect 2792 70514 2912 70530
rect 2780 70508 2912 70514
rect 2832 70502 2912 70508
rect 2964 70508 3016 70514
rect 2780 70450 2832 70456
rect 2964 70450 3016 70456
rect 2700 70378 2820 70394
rect 2700 70372 2832 70378
rect 2700 70366 2780 70372
rect 2780 70314 2832 70320
rect 2582 70204 2890 70224
rect 2582 70202 2588 70204
rect 2644 70202 2668 70204
rect 2724 70202 2748 70204
rect 2804 70202 2828 70204
rect 2884 70202 2890 70204
rect 2644 70150 2646 70202
rect 2826 70150 2828 70202
rect 2582 70148 2588 70150
rect 2644 70148 2668 70150
rect 2724 70148 2748 70150
rect 2804 70148 2828 70150
rect 2884 70148 2890 70150
rect 2582 70128 2890 70148
rect 2872 69964 2924 69970
rect 2872 69906 2924 69912
rect 2884 69306 2912 69906
rect 2976 69426 3004 70450
rect 3068 70310 3096 73902
rect 3160 73846 3188 76230
rect 3252 74118 3280 77590
rect 3344 77042 3372 78367
rect 3896 77330 3924 79183
rect 10138 78704 10194 78713
rect 10138 78639 10194 78648
rect 4066 78024 4122 78033
rect 4066 77959 4122 77968
rect 3974 77616 4030 77625
rect 3974 77551 4030 77560
rect 3988 77518 4016 77551
rect 4080 77518 4108 77959
rect 5845 77820 6153 77840
rect 5845 77818 5851 77820
rect 5907 77818 5931 77820
rect 5987 77818 6011 77820
rect 6067 77818 6091 77820
rect 6147 77818 6153 77820
rect 5907 77766 5909 77818
rect 6089 77766 6091 77818
rect 5845 77764 5851 77766
rect 5907 77764 5931 77766
rect 5987 77764 6011 77766
rect 6067 77764 6091 77766
rect 6147 77764 6153 77766
rect 5845 77744 6153 77764
rect 9109 77820 9417 77840
rect 9109 77818 9115 77820
rect 9171 77818 9195 77820
rect 9251 77818 9275 77820
rect 9331 77818 9355 77820
rect 9411 77818 9417 77820
rect 9171 77766 9173 77818
rect 9353 77766 9355 77818
rect 9109 77764 9115 77766
rect 9171 77764 9195 77766
rect 9251 77764 9275 77766
rect 9331 77764 9355 77766
rect 9411 77764 9417 77766
rect 9109 77744 9417 77764
rect 4712 77648 4764 77654
rect 4712 77590 4764 77596
rect 3976 77512 4028 77518
rect 3976 77454 4028 77460
rect 4068 77512 4120 77518
rect 4068 77454 4120 77460
rect 4620 77376 4672 77382
rect 3896 77302 4108 77330
rect 4620 77318 4672 77324
rect 4080 77058 4108 77302
rect 4213 77276 4521 77296
rect 4213 77274 4219 77276
rect 4275 77274 4299 77276
rect 4355 77274 4379 77276
rect 4435 77274 4459 77276
rect 4515 77274 4521 77276
rect 4275 77222 4277 77274
rect 4457 77222 4459 77274
rect 4213 77220 4219 77222
rect 4275 77220 4299 77222
rect 4355 77220 4379 77222
rect 4435 77220 4459 77222
rect 4515 77220 4521 77222
rect 4213 77200 4521 77220
rect 4080 77042 4200 77058
rect 3332 77036 3384 77042
rect 4080 77036 4212 77042
rect 4080 77030 4160 77036
rect 3332 76978 3384 76984
rect 4160 76978 4212 76984
rect 3424 76900 3476 76906
rect 3424 76842 3476 76848
rect 3332 74860 3384 74866
rect 3332 74802 3384 74808
rect 3344 74254 3372 74802
rect 3332 74248 3384 74254
rect 3332 74190 3384 74196
rect 3240 74112 3292 74118
rect 3240 74054 3292 74060
rect 3148 73840 3200 73846
rect 3148 73782 3200 73788
rect 3240 72072 3292 72078
rect 3240 72014 3292 72020
rect 3252 70394 3280 72014
rect 3344 70514 3372 74190
rect 3436 70650 3464 76842
rect 3516 76832 3568 76838
rect 3516 76774 3568 76780
rect 3976 76832 4028 76838
rect 3976 76774 4028 76780
rect 3528 74934 3556 76774
rect 3884 76560 3936 76566
rect 3884 76502 3936 76508
rect 3608 75948 3660 75954
rect 3608 75890 3660 75896
rect 3516 74928 3568 74934
rect 3516 74870 3568 74876
rect 3620 74361 3648 75890
rect 3792 75200 3844 75206
rect 3792 75142 3844 75148
rect 3606 74352 3662 74361
rect 3606 74287 3662 74296
rect 3804 72146 3832 75142
rect 3896 74866 3924 76502
rect 3988 76498 4016 76774
rect 3976 76492 4028 76498
rect 3976 76434 4028 76440
rect 4213 76188 4521 76208
rect 4213 76186 4219 76188
rect 4275 76186 4299 76188
rect 4355 76186 4379 76188
rect 4435 76186 4459 76188
rect 4515 76186 4521 76188
rect 4275 76134 4277 76186
rect 4457 76134 4459 76186
rect 4213 76132 4219 76134
rect 4275 76132 4299 76134
rect 4355 76132 4379 76134
rect 4435 76132 4459 76134
rect 4515 76132 4521 76134
rect 4213 76112 4521 76132
rect 3976 75336 4028 75342
rect 3976 75278 4028 75284
rect 3988 75041 4016 75278
rect 4213 75100 4521 75120
rect 4213 75098 4219 75100
rect 4275 75098 4299 75100
rect 4355 75098 4379 75100
rect 4435 75098 4459 75100
rect 4515 75098 4521 75100
rect 4275 75046 4277 75098
rect 4457 75046 4459 75098
rect 4213 75044 4219 75046
rect 4275 75044 4299 75046
rect 4355 75044 4379 75046
rect 4435 75044 4459 75046
rect 4515 75044 4521 75046
rect 3974 75032 4030 75041
rect 4213 75024 4521 75044
rect 4632 75002 4660 77318
rect 4724 76090 4752 77590
rect 10152 77518 10180 78639
rect 10966 78024 11022 78033
rect 10966 77959 10968 77968
rect 11020 77959 11022 77968
rect 10968 77930 11020 77936
rect 9404 77512 9456 77518
rect 9404 77454 9456 77460
rect 10140 77512 10192 77518
rect 10140 77454 10192 77460
rect 5080 77376 5132 77382
rect 5080 77318 5132 77324
rect 5092 76634 5120 77318
rect 7477 77276 7785 77296
rect 7477 77274 7483 77276
rect 7539 77274 7563 77276
rect 7619 77274 7643 77276
rect 7699 77274 7723 77276
rect 7779 77274 7785 77276
rect 7539 77222 7541 77274
rect 7721 77222 7723 77274
rect 7477 77220 7483 77222
rect 7539 77220 7563 77222
rect 7619 77220 7643 77222
rect 7699 77220 7723 77222
rect 7779 77220 7785 77222
rect 7477 77200 7785 77220
rect 9416 77217 9444 77454
rect 9402 77208 9458 77217
rect 9402 77143 9458 77152
rect 10140 77036 10192 77042
rect 10140 76978 10192 76984
rect 9864 76832 9916 76838
rect 9864 76774 9916 76780
rect 5845 76732 6153 76752
rect 5845 76730 5851 76732
rect 5907 76730 5931 76732
rect 5987 76730 6011 76732
rect 6067 76730 6091 76732
rect 6147 76730 6153 76732
rect 5907 76678 5909 76730
rect 6089 76678 6091 76730
rect 5845 76676 5851 76678
rect 5907 76676 5931 76678
rect 5987 76676 6011 76678
rect 6067 76676 6091 76678
rect 6147 76676 6153 76678
rect 5845 76656 6153 76676
rect 9109 76732 9417 76752
rect 9109 76730 9115 76732
rect 9171 76730 9195 76732
rect 9251 76730 9275 76732
rect 9331 76730 9355 76732
rect 9411 76730 9417 76732
rect 9171 76678 9173 76730
rect 9353 76678 9355 76730
rect 9109 76676 9115 76678
rect 9171 76676 9195 76678
rect 9251 76676 9275 76678
rect 9331 76676 9355 76678
rect 9411 76676 9417 76678
rect 9109 76656 9417 76676
rect 5080 76628 5132 76634
rect 5080 76570 5132 76576
rect 7477 76188 7785 76208
rect 7477 76186 7483 76188
rect 7539 76186 7563 76188
rect 7619 76186 7643 76188
rect 7699 76186 7723 76188
rect 7779 76186 7785 76188
rect 7539 76134 7541 76186
rect 7721 76134 7723 76186
rect 7477 76132 7483 76134
rect 7539 76132 7563 76134
rect 7619 76132 7643 76134
rect 7699 76132 7723 76134
rect 7779 76132 7785 76134
rect 7477 76112 7785 76132
rect 4712 76084 4764 76090
rect 4712 76026 4764 76032
rect 6368 75948 6420 75954
rect 6368 75890 6420 75896
rect 5845 75644 6153 75664
rect 5845 75642 5851 75644
rect 5907 75642 5931 75644
rect 5987 75642 6011 75644
rect 6067 75642 6091 75644
rect 6147 75642 6153 75644
rect 5907 75590 5909 75642
rect 6089 75590 6091 75642
rect 5845 75588 5851 75590
rect 5907 75588 5931 75590
rect 5987 75588 6011 75590
rect 6067 75588 6091 75590
rect 6147 75588 6153 75590
rect 5845 75568 6153 75588
rect 3974 74967 4030 74976
rect 4620 74996 4672 75002
rect 4620 74938 4672 74944
rect 3884 74860 3936 74866
rect 3884 74802 3936 74808
rect 3792 72140 3844 72146
rect 3792 72082 3844 72088
rect 3424 70644 3476 70650
rect 3424 70586 3476 70592
rect 3332 70508 3384 70514
rect 3332 70450 3384 70456
rect 3516 70508 3568 70514
rect 3516 70450 3568 70456
rect 3148 70372 3200 70378
rect 3252 70366 3372 70394
rect 3148 70314 3200 70320
rect 3056 70304 3108 70310
rect 3056 70246 3108 70252
rect 3068 69970 3096 70246
rect 3056 69964 3108 69970
rect 3056 69906 3108 69912
rect 2964 69420 3016 69426
rect 2964 69362 3016 69368
rect 3160 69358 3188 70314
rect 3240 69896 3292 69902
rect 3240 69838 3292 69844
rect 3252 69426 3280 69838
rect 3344 69562 3372 70366
rect 3528 69873 3556 70450
rect 3608 70304 3660 70310
rect 3608 70246 3660 70252
rect 3514 69864 3570 69873
rect 3514 69799 3570 69808
rect 3516 69760 3568 69766
rect 3516 69702 3568 69708
rect 3332 69556 3384 69562
rect 3332 69498 3384 69504
rect 3240 69420 3292 69426
rect 3240 69362 3292 69368
rect 3148 69352 3200 69358
rect 2884 69278 3004 69306
rect 3148 69294 3200 69300
rect 2582 69116 2890 69136
rect 2582 69114 2588 69116
rect 2644 69114 2668 69116
rect 2724 69114 2748 69116
rect 2804 69114 2828 69116
rect 2884 69114 2890 69116
rect 2644 69062 2646 69114
rect 2826 69062 2828 69114
rect 2582 69060 2588 69062
rect 2644 69060 2668 69062
rect 2724 69060 2748 69062
rect 2804 69060 2828 69062
rect 2884 69060 2890 69062
rect 2582 69040 2890 69060
rect 2976 68882 3004 69278
rect 2964 68876 3016 68882
rect 2964 68818 3016 68824
rect 2964 68740 3016 68746
rect 2964 68682 3016 68688
rect 2582 68028 2890 68048
rect 2582 68026 2588 68028
rect 2644 68026 2668 68028
rect 2724 68026 2748 68028
rect 2804 68026 2828 68028
rect 2884 68026 2890 68028
rect 2644 67974 2646 68026
rect 2826 67974 2828 68026
rect 2582 67972 2588 67974
rect 2644 67972 2668 67974
rect 2724 67972 2748 67974
rect 2804 67972 2828 67974
rect 2884 67972 2890 67974
rect 2582 67952 2890 67972
rect 2976 67658 3004 68682
rect 3160 67862 3188 69294
rect 3240 68468 3292 68474
rect 3240 68410 3292 68416
rect 3148 67856 3200 67862
rect 3148 67798 3200 67804
rect 2964 67652 3016 67658
rect 2964 67594 3016 67600
rect 3056 67652 3108 67658
rect 3056 67594 3108 67600
rect 2976 67250 3004 67594
rect 2964 67244 3016 67250
rect 2964 67186 3016 67192
rect 2582 66940 2890 66960
rect 2582 66938 2588 66940
rect 2644 66938 2668 66940
rect 2724 66938 2748 66940
rect 2804 66938 2828 66940
rect 2884 66938 2890 66940
rect 2644 66886 2646 66938
rect 2826 66886 2828 66938
rect 2582 66884 2588 66886
rect 2644 66884 2668 66886
rect 2724 66884 2748 66886
rect 2804 66884 2828 66886
rect 2884 66884 2890 66886
rect 2582 66864 2890 66884
rect 2962 66736 3018 66745
rect 2962 66671 3018 66680
rect 2976 66638 3004 66671
rect 2964 66632 3016 66638
rect 2964 66574 3016 66580
rect 3068 66178 3096 67594
rect 3148 67244 3200 67250
rect 3148 67186 3200 67192
rect 2976 66150 3096 66178
rect 2582 65852 2890 65872
rect 2582 65850 2588 65852
rect 2644 65850 2668 65852
rect 2724 65850 2748 65852
rect 2804 65850 2828 65852
rect 2884 65850 2890 65852
rect 2644 65798 2646 65850
rect 2826 65798 2828 65850
rect 2582 65796 2588 65798
rect 2644 65796 2668 65798
rect 2724 65796 2748 65798
rect 2804 65796 2828 65798
rect 2884 65796 2890 65798
rect 2582 65776 2890 65796
rect 2582 64764 2890 64784
rect 2582 64762 2588 64764
rect 2644 64762 2668 64764
rect 2724 64762 2748 64764
rect 2804 64762 2828 64764
rect 2884 64762 2890 64764
rect 2644 64710 2646 64762
rect 2826 64710 2828 64762
rect 2582 64708 2588 64710
rect 2644 64708 2668 64710
rect 2724 64708 2748 64710
rect 2804 64708 2828 64710
rect 2884 64708 2890 64710
rect 2582 64688 2890 64708
rect 2582 63676 2890 63696
rect 2582 63674 2588 63676
rect 2644 63674 2668 63676
rect 2724 63674 2748 63676
rect 2804 63674 2828 63676
rect 2884 63674 2890 63676
rect 2644 63622 2646 63674
rect 2826 63622 2828 63674
rect 2582 63620 2588 63622
rect 2644 63620 2668 63622
rect 2724 63620 2748 63622
rect 2804 63620 2828 63622
rect 2884 63620 2890 63622
rect 2582 63600 2890 63620
rect 2870 63472 2926 63481
rect 2870 63407 2872 63416
rect 2924 63407 2926 63416
rect 2872 63378 2924 63384
rect 2872 63300 2924 63306
rect 2872 63242 2924 63248
rect 2884 63209 2912 63242
rect 2870 63200 2926 63209
rect 2870 63135 2926 63144
rect 2582 62588 2890 62608
rect 2582 62586 2588 62588
rect 2644 62586 2668 62588
rect 2724 62586 2748 62588
rect 2804 62586 2828 62588
rect 2884 62586 2890 62588
rect 2644 62534 2646 62586
rect 2826 62534 2828 62586
rect 2582 62532 2588 62534
rect 2644 62532 2668 62534
rect 2724 62532 2748 62534
rect 2804 62532 2828 62534
rect 2884 62532 2890 62534
rect 2582 62512 2890 62532
rect 2976 61878 3004 66150
rect 3056 65408 3108 65414
rect 3056 65350 3108 65356
rect 3068 65113 3096 65350
rect 3054 65104 3110 65113
rect 3054 65039 3110 65048
rect 3056 65000 3108 65006
rect 3160 64954 3188 67186
rect 3108 64948 3188 64954
rect 3056 64942 3188 64948
rect 3068 64926 3188 64942
rect 3068 62830 3096 64926
rect 3148 63776 3200 63782
rect 3148 63718 3200 63724
rect 3160 63345 3188 63718
rect 3146 63336 3202 63345
rect 3146 63271 3202 63280
rect 3056 62824 3108 62830
rect 3056 62766 3108 62772
rect 3056 62688 3108 62694
rect 3056 62630 3108 62636
rect 2964 61872 3016 61878
rect 2964 61814 3016 61820
rect 2964 61600 3016 61606
rect 2964 61542 3016 61548
rect 2582 61500 2890 61520
rect 2582 61498 2588 61500
rect 2644 61498 2668 61500
rect 2724 61498 2748 61500
rect 2804 61498 2828 61500
rect 2884 61498 2890 61500
rect 2644 61446 2646 61498
rect 2826 61446 2828 61498
rect 2582 61444 2588 61446
rect 2644 61444 2668 61446
rect 2724 61444 2748 61446
rect 2804 61444 2828 61446
rect 2884 61444 2890 61446
rect 2582 61424 2890 61444
rect 2780 61056 2832 61062
rect 2780 60998 2832 61004
rect 2792 60625 2820 60998
rect 2976 60761 3004 61542
rect 2962 60752 3018 60761
rect 2962 60687 3018 60696
rect 2778 60616 2834 60625
rect 2778 60551 2834 60560
rect 2582 60412 2890 60432
rect 2582 60410 2588 60412
rect 2644 60410 2668 60412
rect 2724 60410 2748 60412
rect 2804 60410 2828 60412
rect 2884 60410 2890 60412
rect 2644 60358 2646 60410
rect 2826 60358 2828 60410
rect 2582 60356 2588 60358
rect 2644 60356 2668 60358
rect 2724 60356 2748 60358
rect 2804 60356 2828 60358
rect 2884 60356 2890 60358
rect 2582 60336 2890 60356
rect 2964 60036 3016 60042
rect 2964 59978 3016 59984
rect 2872 59968 2924 59974
rect 2872 59910 2924 59916
rect 2516 59758 2636 59786
rect 2884 59770 2912 59910
rect 2608 59514 2636 59758
rect 2872 59764 2924 59770
rect 2872 59706 2924 59712
rect 2516 59486 2636 59514
rect 2412 57588 2464 57594
rect 2412 57530 2464 57536
rect 2320 57452 2372 57458
rect 2320 57394 2372 57400
rect 2332 56982 2360 57394
rect 2320 56976 2372 56982
rect 2320 56918 2372 56924
rect 2516 56778 2544 59486
rect 2582 59324 2890 59344
rect 2582 59322 2588 59324
rect 2644 59322 2668 59324
rect 2724 59322 2748 59324
rect 2804 59322 2828 59324
rect 2884 59322 2890 59324
rect 2644 59270 2646 59322
rect 2826 59270 2828 59322
rect 2582 59268 2588 59270
rect 2644 59268 2668 59270
rect 2724 59268 2748 59270
rect 2804 59268 2828 59270
rect 2884 59268 2890 59270
rect 2582 59248 2890 59268
rect 2582 58236 2890 58256
rect 2582 58234 2588 58236
rect 2644 58234 2668 58236
rect 2724 58234 2748 58236
rect 2804 58234 2828 58236
rect 2884 58234 2890 58236
rect 2644 58182 2646 58234
rect 2826 58182 2828 58234
rect 2582 58180 2588 58182
rect 2644 58180 2668 58182
rect 2724 58180 2748 58182
rect 2804 58180 2828 58182
rect 2884 58180 2890 58182
rect 2582 58160 2890 58180
rect 2872 58064 2924 58070
rect 2872 58006 2924 58012
rect 2780 57792 2832 57798
rect 2778 57760 2780 57769
rect 2832 57760 2834 57769
rect 2778 57695 2834 57704
rect 2884 57361 2912 58006
rect 2870 57352 2926 57361
rect 2870 57287 2926 57296
rect 2582 57148 2890 57168
rect 2582 57146 2588 57148
rect 2644 57146 2668 57148
rect 2724 57146 2748 57148
rect 2804 57146 2828 57148
rect 2884 57146 2890 57148
rect 2644 57094 2646 57146
rect 2826 57094 2828 57146
rect 2582 57092 2588 57094
rect 2644 57092 2668 57094
rect 2724 57092 2748 57094
rect 2804 57092 2828 57094
rect 2884 57092 2890 57094
rect 2582 57072 2890 57092
rect 2780 56976 2832 56982
rect 2780 56918 2832 56924
rect 2596 56908 2648 56914
rect 2596 56850 2648 56856
rect 2608 56794 2636 56850
rect 2792 56794 2820 56918
rect 2504 56772 2556 56778
rect 2608 56766 2820 56794
rect 2504 56714 2556 56720
rect 2976 56658 3004 59978
rect 2792 56630 3004 56658
rect 2792 56438 2820 56630
rect 3068 56488 3096 62630
rect 3148 61872 3200 61878
rect 3148 61814 3200 61820
rect 3160 60042 3188 61814
rect 3148 60036 3200 60042
rect 3148 59978 3200 59984
rect 3148 59764 3200 59770
rect 3148 59706 3200 59712
rect 2884 56460 3096 56488
rect 2320 56432 2372 56438
rect 2320 56374 2372 56380
rect 2780 56432 2832 56438
rect 2780 56374 2832 56380
rect 2226 54632 2282 54641
rect 2226 54567 2282 54576
rect 2228 54528 2280 54534
rect 2228 54470 2280 54476
rect 2240 54369 2268 54470
rect 2226 54360 2282 54369
rect 2226 54295 2282 54304
rect 2136 53440 2188 53446
rect 2136 53382 2188 53388
rect 2332 52986 2360 56374
rect 2884 56234 2912 56460
rect 3160 56273 3188 59706
rect 3252 57497 3280 68410
rect 3344 68338 3372 69498
rect 3332 68332 3384 68338
rect 3332 68274 3384 68280
rect 3424 68332 3476 68338
rect 3424 68274 3476 68280
rect 3344 67386 3372 68274
rect 3436 68241 3464 68274
rect 3422 68232 3478 68241
rect 3422 68167 3478 68176
rect 3424 67856 3476 67862
rect 3424 67798 3476 67804
rect 3332 67380 3384 67386
rect 3332 67322 3384 67328
rect 3332 66632 3384 66638
rect 3332 66574 3384 66580
rect 3344 60858 3372 66574
rect 3436 64394 3464 67798
rect 3424 64388 3476 64394
rect 3424 64330 3476 64336
rect 3436 62098 3464 64330
rect 3528 62218 3556 69702
rect 3620 66638 3648 70246
rect 3700 69760 3752 69766
rect 3700 69702 3752 69708
rect 3608 66632 3660 66638
rect 3608 66574 3660 66580
rect 3608 66496 3660 66502
rect 3608 66438 3660 66444
rect 3516 62212 3568 62218
rect 3516 62154 3568 62160
rect 3436 62070 3556 62098
rect 3424 61192 3476 61198
rect 3424 61134 3476 61140
rect 3332 60852 3384 60858
rect 3332 60794 3384 60800
rect 3330 60752 3386 60761
rect 3330 60687 3386 60696
rect 3344 60654 3372 60687
rect 3332 60648 3384 60654
rect 3332 60590 3384 60596
rect 3238 57488 3294 57497
rect 3344 57458 3372 60590
rect 3238 57423 3294 57432
rect 3332 57452 3384 57458
rect 3332 57394 3384 57400
rect 3344 56982 3372 57394
rect 3332 56976 3384 56982
rect 3332 56918 3384 56924
rect 3240 56296 3292 56302
rect 3146 56264 3202 56273
rect 2872 56228 2924 56234
rect 2872 56170 2924 56176
rect 3056 56228 3108 56234
rect 3240 56238 3292 56244
rect 3146 56199 3202 56208
rect 3056 56170 3108 56176
rect 2582 56060 2890 56080
rect 2582 56058 2588 56060
rect 2644 56058 2668 56060
rect 2724 56058 2748 56060
rect 2804 56058 2828 56060
rect 2884 56058 2890 56060
rect 2644 56006 2646 56058
rect 2826 56006 2828 56058
rect 2582 56004 2588 56006
rect 2644 56004 2668 56006
rect 2724 56004 2748 56006
rect 2804 56004 2828 56006
rect 2884 56004 2890 56006
rect 2582 55984 2890 56004
rect 2412 55956 2464 55962
rect 2412 55898 2464 55904
rect 2148 52958 2360 52986
rect 2148 51882 2176 52958
rect 2228 52896 2280 52902
rect 2228 52838 2280 52844
rect 2240 52601 2268 52838
rect 2424 52698 2452 55898
rect 2504 55616 2556 55622
rect 2504 55558 2556 55564
rect 2780 55616 2832 55622
rect 2780 55558 2832 55564
rect 2516 54194 2544 55558
rect 2792 55350 2820 55558
rect 2780 55344 2832 55350
rect 2780 55286 2832 55292
rect 2778 55176 2834 55185
rect 2778 55111 2780 55120
rect 2832 55111 2834 55120
rect 2780 55082 2832 55088
rect 2582 54972 2890 54992
rect 2582 54970 2588 54972
rect 2644 54970 2668 54972
rect 2724 54970 2748 54972
rect 2804 54970 2828 54972
rect 2884 54970 2890 54972
rect 2644 54918 2646 54970
rect 2826 54918 2828 54970
rect 2582 54916 2588 54918
rect 2644 54916 2668 54918
rect 2724 54916 2748 54918
rect 2804 54916 2828 54918
rect 2884 54916 2890 54918
rect 2582 54896 2890 54916
rect 3068 54330 3096 56170
rect 3148 56160 3200 56166
rect 3148 56102 3200 56108
rect 3160 55865 3188 56102
rect 3146 55856 3202 55865
rect 3146 55791 3202 55800
rect 3148 55684 3200 55690
rect 3148 55626 3200 55632
rect 3160 55457 3188 55626
rect 3146 55448 3202 55457
rect 3146 55383 3202 55392
rect 3252 55350 3280 56238
rect 3344 55894 3372 56918
rect 3332 55888 3384 55894
rect 3332 55830 3384 55836
rect 3240 55344 3292 55350
rect 3240 55286 3292 55292
rect 3056 54324 3108 54330
rect 3056 54266 3108 54272
rect 2504 54188 2556 54194
rect 2504 54130 2556 54136
rect 2964 54188 3016 54194
rect 2964 54130 3016 54136
rect 3332 54188 3384 54194
rect 3332 54130 3384 54136
rect 2582 53884 2890 53904
rect 2582 53882 2588 53884
rect 2644 53882 2668 53884
rect 2724 53882 2748 53884
rect 2804 53882 2828 53884
rect 2884 53882 2890 53884
rect 2644 53830 2646 53882
rect 2826 53830 2828 53882
rect 2582 53828 2588 53830
rect 2644 53828 2668 53830
rect 2724 53828 2748 53830
rect 2804 53828 2828 53830
rect 2884 53828 2890 53830
rect 2582 53808 2890 53828
rect 2778 53544 2834 53553
rect 2778 53479 2834 53488
rect 2792 53446 2820 53479
rect 2780 53440 2832 53446
rect 2780 53382 2832 53388
rect 2504 53236 2556 53242
rect 2504 53178 2556 53184
rect 2412 52692 2464 52698
rect 2412 52634 2464 52640
rect 2226 52592 2282 52601
rect 2226 52527 2282 52536
rect 2228 52488 2280 52494
rect 2228 52430 2280 52436
rect 2412 52488 2464 52494
rect 2412 52430 2464 52436
rect 2136 51876 2188 51882
rect 2136 51818 2188 51824
rect 2240 51456 2268 52430
rect 2320 52352 2372 52358
rect 2320 52294 2372 52300
rect 2332 52018 2360 52294
rect 2320 52012 2372 52018
rect 2320 51954 2372 51960
rect 2320 51876 2372 51882
rect 2320 51818 2372 51824
rect 2148 51428 2268 51456
rect 2148 51241 2176 51428
rect 2226 51368 2282 51377
rect 2226 51303 2282 51312
rect 2240 51270 2268 51303
rect 2228 51264 2280 51270
rect 2134 51232 2190 51241
rect 2228 51206 2280 51212
rect 2134 51167 2190 51176
rect 2228 51060 2280 51066
rect 1964 51020 2228 51048
rect 2228 51002 2280 51008
rect 2226 50960 2282 50969
rect 2226 50895 2228 50904
rect 2280 50895 2282 50904
rect 2228 50866 2280 50872
rect 2134 50824 2190 50833
rect 1952 50788 2004 50794
rect 2134 50759 2190 50768
rect 1952 50730 2004 50736
rect 1860 50312 1912 50318
rect 1860 50254 1912 50260
rect 1768 49972 1820 49978
rect 1768 49914 1820 49920
rect 1964 49858 1992 50730
rect 2042 50688 2098 50697
rect 2042 50623 2098 50632
rect 1872 49830 1992 49858
rect 1676 49768 1728 49774
rect 1728 49716 1808 49722
rect 1676 49710 1808 49716
rect 1688 49694 1808 49710
rect 1596 49558 1716 49586
rect 1584 49428 1636 49434
rect 1584 49370 1636 49376
rect 1400 49224 1452 49230
rect 1400 49166 1452 49172
rect 1400 49088 1452 49094
rect 1400 49030 1452 49036
rect 1412 43790 1440 49030
rect 1492 48544 1544 48550
rect 1492 48486 1544 48492
rect 1504 48385 1532 48486
rect 1490 48376 1546 48385
rect 1490 48311 1546 48320
rect 1492 48000 1544 48006
rect 1492 47942 1544 47948
rect 1504 47841 1532 47942
rect 1490 47832 1546 47841
rect 1490 47767 1546 47776
rect 1492 47456 1544 47462
rect 1492 47398 1544 47404
rect 1504 47025 1532 47398
rect 1490 47016 1546 47025
rect 1490 46951 1546 46960
rect 1492 46912 1544 46918
rect 1492 46854 1544 46860
rect 1504 46617 1532 46854
rect 1490 46608 1546 46617
rect 1490 46543 1546 46552
rect 1492 46368 1544 46374
rect 1492 46310 1544 46316
rect 1504 46209 1532 46310
rect 1490 46200 1546 46209
rect 1490 46135 1546 46144
rect 1492 45280 1544 45286
rect 1490 45248 1492 45257
rect 1544 45248 1546 45257
rect 1490 45183 1546 45192
rect 1596 44520 1624 49370
rect 1504 44492 1624 44520
rect 1400 43784 1452 43790
rect 1400 43726 1452 43732
rect 1320 43608 1440 43636
rect 1412 42650 1440 43608
rect 1504 43246 1532 44492
rect 1582 44432 1638 44441
rect 1582 44367 1638 44376
rect 1596 43994 1624 44367
rect 1584 43988 1636 43994
rect 1584 43930 1636 43936
rect 1492 43240 1544 43246
rect 1492 43182 1544 43188
rect 1492 43104 1544 43110
rect 1492 43046 1544 43052
rect 1320 42622 1440 42650
rect 1320 41818 1348 42622
rect 1400 42560 1452 42566
rect 1400 42502 1452 42508
rect 1412 41857 1440 42502
rect 1504 42265 1532 43046
rect 1490 42256 1546 42265
rect 1490 42191 1546 42200
rect 1492 42016 1544 42022
rect 1492 41958 1544 41964
rect 1398 41848 1454 41857
rect 1308 41812 1360 41818
rect 1398 41783 1454 41792
rect 1308 41754 1360 41760
rect 1400 41472 1452 41478
rect 1504 41449 1532 41958
rect 1400 41414 1452 41420
rect 1490 41440 1546 41449
rect 1412 40633 1440 41414
rect 1490 41375 1546 41384
rect 1688 41274 1716 49558
rect 1780 49434 1808 49694
rect 1768 49428 1820 49434
rect 1768 49370 1820 49376
rect 1768 48068 1820 48074
rect 1768 48010 1820 48016
rect 1780 45966 1808 48010
rect 1872 46322 1900 49830
rect 1952 49428 2004 49434
rect 1952 49370 2004 49376
rect 1964 49230 1992 49370
rect 1952 49224 2004 49230
rect 1952 49166 2004 49172
rect 1950 49056 2006 49065
rect 1950 48991 2006 49000
rect 1964 48822 1992 48991
rect 1952 48816 2004 48822
rect 1952 48758 2004 48764
rect 2056 48226 2084 50623
rect 1964 48198 2084 48226
rect 1964 46714 1992 48198
rect 2044 48136 2096 48142
rect 2044 48078 2096 48084
rect 2056 47734 2084 48078
rect 2044 47728 2096 47734
rect 2044 47670 2096 47676
rect 1952 46708 2004 46714
rect 1952 46650 2004 46656
rect 1872 46294 2084 46322
rect 1860 46164 1912 46170
rect 1860 46106 1912 46112
rect 1768 45960 1820 45966
rect 1768 45902 1820 45908
rect 1780 44878 1808 45902
rect 1768 44872 1820 44878
rect 1768 44814 1820 44820
rect 1780 44402 1808 44814
rect 1768 44396 1820 44402
rect 1768 44338 1820 44344
rect 1768 43716 1820 43722
rect 1768 43658 1820 43664
rect 1780 43314 1808 43658
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1768 43172 1820 43178
rect 1768 43114 1820 43120
rect 1780 42106 1808 43114
rect 1872 42265 1900 46106
rect 1952 45824 2004 45830
rect 1952 45766 2004 45772
rect 1858 42256 1914 42265
rect 1964 42242 1992 45766
rect 2056 45121 2084 46294
rect 2148 46170 2176 50759
rect 2228 50312 2280 50318
rect 2228 50254 2280 50260
rect 2240 49842 2268 50254
rect 2228 49836 2280 49842
rect 2228 49778 2280 49784
rect 2240 49366 2268 49778
rect 2228 49360 2280 49366
rect 2228 49302 2280 49308
rect 2226 49192 2282 49201
rect 2226 49127 2282 49136
rect 2240 48890 2268 49127
rect 2228 48884 2280 48890
rect 2228 48826 2280 48832
rect 2228 48748 2280 48754
rect 2228 48690 2280 48696
rect 2240 48657 2268 48690
rect 2226 48648 2282 48657
rect 2226 48583 2282 48592
rect 2228 47456 2280 47462
rect 2226 47424 2228 47433
rect 2280 47424 2282 47433
rect 2226 47359 2282 47368
rect 2332 47258 2360 51818
rect 2424 51542 2452 52430
rect 2412 51536 2464 51542
rect 2412 51478 2464 51484
rect 2516 51320 2544 53178
rect 2582 52796 2890 52816
rect 2582 52794 2588 52796
rect 2644 52794 2668 52796
rect 2724 52794 2748 52796
rect 2804 52794 2828 52796
rect 2884 52794 2890 52796
rect 2644 52742 2646 52794
rect 2826 52742 2828 52794
rect 2582 52740 2588 52742
rect 2644 52740 2668 52742
rect 2724 52740 2748 52742
rect 2804 52740 2828 52742
rect 2884 52740 2890 52742
rect 2582 52720 2890 52740
rect 2872 52420 2924 52426
rect 2976 52408 3004 54130
rect 3054 53000 3110 53009
rect 3054 52935 3056 52944
rect 3108 52935 3110 52944
rect 3056 52906 3108 52912
rect 3056 52488 3108 52494
rect 3056 52430 3108 52436
rect 2924 52380 3004 52408
rect 2872 52362 2924 52368
rect 2884 51882 2912 52362
rect 3068 52018 3096 52430
rect 3148 52420 3200 52426
rect 3148 52362 3200 52368
rect 3160 52154 3188 52362
rect 3148 52148 3200 52154
rect 3148 52090 3200 52096
rect 2964 52012 3016 52018
rect 2964 51954 3016 51960
rect 3056 52012 3108 52018
rect 3056 51954 3108 51960
rect 2872 51876 2924 51882
rect 2872 51818 2924 51824
rect 2582 51708 2890 51728
rect 2582 51706 2588 51708
rect 2644 51706 2668 51708
rect 2724 51706 2748 51708
rect 2804 51706 2828 51708
rect 2884 51706 2890 51708
rect 2644 51654 2646 51706
rect 2826 51654 2828 51706
rect 2582 51652 2588 51654
rect 2644 51652 2668 51654
rect 2724 51652 2748 51654
rect 2804 51652 2828 51654
rect 2884 51652 2890 51654
rect 2582 51632 2890 51652
rect 2688 51536 2740 51542
rect 2976 51524 3004 51954
rect 3148 51876 3200 51882
rect 3148 51818 3200 51824
rect 2688 51478 2740 51484
rect 2884 51496 3004 51524
rect 2424 51292 2544 51320
rect 2424 50454 2452 51292
rect 2502 51096 2558 51105
rect 2502 51031 2558 51040
rect 2516 50930 2544 51031
rect 2504 50924 2556 50930
rect 2504 50866 2556 50872
rect 2502 50824 2558 50833
rect 2700 50794 2728 51478
rect 2780 51400 2832 51406
rect 2780 51342 2832 51348
rect 2792 50969 2820 51342
rect 2778 50960 2834 50969
rect 2778 50895 2780 50904
rect 2832 50895 2834 50904
rect 2780 50866 2832 50872
rect 2792 50835 2820 50866
rect 2884 50833 2912 51496
rect 3160 51474 3188 51818
rect 3148 51468 3200 51474
rect 3148 51410 3200 51416
rect 3056 51400 3108 51406
rect 3056 51342 3108 51348
rect 2964 51332 3016 51338
rect 2964 51274 3016 51280
rect 2870 50824 2926 50833
rect 2502 50759 2558 50768
rect 2688 50788 2740 50794
rect 2412 50448 2464 50454
rect 2412 50390 2464 50396
rect 2412 49836 2464 49842
rect 2412 49778 2464 49784
rect 2424 49745 2452 49778
rect 2410 49736 2466 49745
rect 2410 49671 2466 49680
rect 2412 49632 2464 49638
rect 2410 49600 2412 49609
rect 2464 49600 2466 49609
rect 2410 49535 2466 49544
rect 2412 48340 2464 48346
rect 2412 48282 2464 48288
rect 2320 47252 2372 47258
rect 2320 47194 2372 47200
rect 2424 47138 2452 48282
rect 2240 47110 2452 47138
rect 2136 46164 2188 46170
rect 2136 46106 2188 46112
rect 2134 46064 2190 46073
rect 2134 45999 2190 46008
rect 2148 45966 2176 45999
rect 2136 45960 2188 45966
rect 2136 45902 2188 45908
rect 2042 45112 2098 45121
rect 2042 45047 2098 45056
rect 2044 44940 2096 44946
rect 2044 44882 2096 44888
rect 2056 42378 2084 44882
rect 2148 42906 2176 45902
rect 2240 43790 2268 47110
rect 2320 47048 2372 47054
rect 2320 46990 2372 46996
rect 2332 46481 2360 46990
rect 2412 46708 2464 46714
rect 2412 46650 2464 46656
rect 2318 46472 2374 46481
rect 2318 46407 2374 46416
rect 2320 45960 2372 45966
rect 2320 45902 2372 45908
rect 2228 43784 2280 43790
rect 2228 43726 2280 43732
rect 2228 43648 2280 43654
rect 2332 43636 2360 45902
rect 2424 45830 2452 46650
rect 2412 45824 2464 45830
rect 2412 45766 2464 45772
rect 2410 45656 2466 45665
rect 2410 45591 2466 45600
rect 2424 44946 2452 45591
rect 2412 44940 2464 44946
rect 2412 44882 2464 44888
rect 2410 44840 2466 44849
rect 2410 44775 2466 44784
rect 2424 44742 2452 44775
rect 2412 44736 2464 44742
rect 2412 44678 2464 44684
rect 2412 44192 2464 44198
rect 2412 44134 2464 44140
rect 2424 44033 2452 44134
rect 2410 44024 2466 44033
rect 2410 43959 2466 43968
rect 2332 43608 2452 43636
rect 2228 43590 2280 43596
rect 2240 43217 2268 43590
rect 2318 43480 2374 43489
rect 2318 43415 2374 43424
rect 2226 43208 2282 43217
rect 2226 43143 2282 43152
rect 2136 42900 2188 42906
rect 2136 42842 2188 42848
rect 2332 42702 2360 43415
rect 2320 42696 2372 42702
rect 2226 42664 2282 42673
rect 2320 42638 2372 42644
rect 2226 42599 2282 42608
rect 2240 42566 2268 42599
rect 2228 42560 2280 42566
rect 2228 42502 2280 42508
rect 2056 42350 2360 42378
rect 1964 42214 2268 42242
rect 1858 42191 1914 42200
rect 2042 42120 2098 42129
rect 1780 42078 1992 42106
rect 1858 41848 1914 41857
rect 1858 41783 1914 41792
rect 1768 41608 1820 41614
rect 1768 41550 1820 41556
rect 1780 41313 1808 41550
rect 1766 41304 1822 41313
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1676 41268 1728 41274
rect 1766 41239 1822 41248
rect 1676 41210 1728 41216
rect 1492 41132 1544 41138
rect 1492 41074 1544 41080
rect 1398 40624 1454 40633
rect 1398 40559 1454 40568
rect 1504 40474 1532 41074
rect 1412 40446 1532 40474
rect 1412 39386 1440 40446
rect 1492 40384 1544 40390
rect 1492 40326 1544 40332
rect 1320 39358 1440 39386
rect 1320 37890 1348 39358
rect 1400 39296 1452 39302
rect 1504 39273 1532 40326
rect 1400 39238 1452 39244
rect 1490 39264 1546 39273
rect 1412 38049 1440 39238
rect 1490 39199 1546 39208
rect 1398 38040 1454 38049
rect 1398 37975 1454 37984
rect 1320 37862 1440 37890
rect 1412 36938 1440 37862
rect 1492 37664 1544 37670
rect 1492 37606 1544 37612
rect 1504 37097 1532 37606
rect 1596 37262 1624 41210
rect 1674 41168 1730 41177
rect 1674 41103 1730 41112
rect 1768 41132 1820 41138
rect 1688 40526 1716 41103
rect 1768 41074 1820 41080
rect 1676 40520 1728 40526
rect 1676 40462 1728 40468
rect 1676 40384 1728 40390
rect 1676 40326 1728 40332
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 1688 37210 1716 40326
rect 1780 38010 1808 41074
rect 1872 40390 1900 41783
rect 1860 40384 1912 40390
rect 1860 40326 1912 40332
rect 1860 40044 1912 40050
rect 1860 39986 1912 39992
rect 1872 39370 1900 39986
rect 1860 39364 1912 39370
rect 1860 39306 1912 39312
rect 1872 38962 1900 39306
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 1860 38820 1912 38826
rect 1860 38762 1912 38768
rect 1768 38004 1820 38010
rect 1768 37946 1820 37952
rect 1490 37088 1546 37097
rect 1490 37023 1546 37032
rect 1412 36910 1532 36938
rect 1400 36576 1452 36582
rect 1400 36518 1452 36524
rect 1412 35873 1440 36518
rect 1504 36145 1532 36910
rect 1490 36136 1546 36145
rect 1490 36071 1546 36080
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1398 35864 1454 35873
rect 1398 35799 1454 35808
rect 1398 35728 1454 35737
rect 1398 35663 1454 35672
rect 1412 33402 1440 35663
rect 1504 35465 1532 35974
rect 1490 35456 1546 35465
rect 1490 35391 1546 35400
rect 1490 35048 1546 35057
rect 1490 34983 1546 34992
rect 1504 34950 1532 34983
rect 1492 34944 1544 34950
rect 1492 34886 1544 34892
rect 1596 34746 1624 37198
rect 1688 37182 1808 37210
rect 1676 37120 1728 37126
rect 1676 37062 1728 37068
rect 1688 36922 1716 37062
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 1780 35698 1808 37182
rect 1768 35692 1820 35698
rect 1688 35652 1768 35680
rect 1584 34740 1636 34746
rect 1584 34682 1636 34688
rect 1584 34604 1636 34610
rect 1584 34546 1636 34552
rect 1492 33856 1544 33862
rect 1492 33798 1544 33804
rect 1320 33374 1440 33402
rect 1216 32904 1268 32910
rect 1216 32846 1268 32852
rect 1216 32768 1268 32774
rect 1216 32710 1268 32716
rect 1228 31929 1256 32710
rect 1320 32570 1348 33374
rect 1400 33312 1452 33318
rect 1504 33289 1532 33798
rect 1400 33254 1452 33260
rect 1490 33280 1546 33289
rect 1308 32564 1360 32570
rect 1308 32506 1360 32512
rect 1412 32473 1440 33254
rect 1490 33215 1546 33224
rect 1398 32464 1454 32473
rect 1308 32428 1360 32434
rect 1398 32399 1454 32408
rect 1308 32370 1360 32376
rect 1214 31920 1270 31929
rect 1214 31855 1270 31864
rect 1216 26376 1268 26382
rect 1216 26318 1268 26324
rect 1124 25492 1176 25498
rect 1124 25434 1176 25440
rect 1228 24313 1256 26318
rect 1214 24304 1270 24313
rect 1214 24239 1270 24248
rect 1032 23792 1084 23798
rect 1032 23734 1084 23740
rect 1216 23724 1268 23730
rect 1216 23666 1268 23672
rect 1228 22137 1256 23666
rect 1214 22128 1270 22137
rect 1214 22063 1270 22072
rect 1216 17196 1268 17202
rect 1216 17138 1268 17144
rect 1124 16584 1176 16590
rect 1124 16526 1176 16532
rect 1136 14793 1164 16526
rect 1228 15609 1256 17138
rect 1214 15600 1270 15609
rect 1214 15535 1270 15544
rect 1122 14784 1178 14793
rect 1122 14719 1178 14728
rect 1320 11778 1348 32370
rect 1596 32314 1624 34546
rect 1412 32286 1624 32314
rect 1412 30054 1440 32286
rect 1492 32224 1544 32230
rect 1688 32178 1716 35652
rect 1768 35634 1820 35640
rect 1768 34196 1820 34202
rect 1768 34138 1820 34144
rect 1492 32166 1544 32172
rect 1504 32026 1532 32166
rect 1596 32150 1716 32178
rect 1492 32020 1544 32026
rect 1492 31962 1544 31968
rect 1490 30696 1546 30705
rect 1490 30631 1546 30640
rect 1504 30598 1532 30631
rect 1492 30592 1544 30598
rect 1492 30534 1544 30540
rect 1492 30388 1544 30394
rect 1492 30330 1544 30336
rect 1400 30048 1452 30054
rect 1400 29990 1452 29996
rect 1400 28960 1452 28966
rect 1400 28902 1452 28908
rect 1412 28121 1440 28902
rect 1504 28150 1532 30330
rect 1596 29850 1624 32150
rect 1674 32056 1730 32065
rect 1674 31991 1730 32000
rect 1688 30394 1716 31991
rect 1780 31793 1808 34138
rect 1766 31784 1822 31793
rect 1766 31719 1822 31728
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 1676 30388 1728 30394
rect 1676 30330 1728 30336
rect 1676 30252 1728 30258
rect 1676 30194 1728 30200
rect 1688 29850 1716 30194
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1676 29844 1728 29850
rect 1676 29786 1728 29792
rect 1584 29708 1636 29714
rect 1584 29650 1636 29656
rect 1492 28144 1544 28150
rect 1398 28112 1454 28121
rect 1492 28086 1544 28092
rect 1398 28047 1454 28056
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 25945 1440 27406
rect 1596 26450 1624 29650
rect 1780 29646 1808 30534
rect 1872 30326 1900 38762
rect 1964 33998 1992 42078
rect 2042 42055 2098 42064
rect 1952 33992 2004 33998
rect 1952 33934 2004 33940
rect 1952 33516 2004 33522
rect 1952 33458 2004 33464
rect 1964 32502 1992 33458
rect 2056 32910 2084 42055
rect 2134 41304 2190 41313
rect 2134 41239 2190 41248
rect 2148 38298 2176 41239
rect 2240 41206 2268 42214
rect 2332 41313 2360 42350
rect 2318 41304 2374 41313
rect 2318 41239 2374 41248
rect 2228 41200 2280 41206
rect 2228 41142 2280 41148
rect 2318 41032 2374 41041
rect 2318 40967 2320 40976
rect 2372 40967 2374 40976
rect 2320 40938 2372 40944
rect 2320 40384 2372 40390
rect 2320 40326 2372 40332
rect 2332 39681 2360 40326
rect 2318 39672 2374 39681
rect 2318 39607 2374 39616
rect 2424 39522 2452 43608
rect 2516 41414 2544 50759
rect 2870 50759 2926 50768
rect 2688 50730 2740 50736
rect 2582 50620 2890 50640
rect 2582 50618 2588 50620
rect 2644 50618 2668 50620
rect 2724 50618 2748 50620
rect 2804 50618 2828 50620
rect 2884 50618 2890 50620
rect 2644 50566 2646 50618
rect 2826 50566 2828 50618
rect 2582 50564 2588 50566
rect 2644 50564 2668 50566
rect 2724 50564 2748 50566
rect 2804 50564 2828 50566
rect 2884 50564 2890 50566
rect 2582 50544 2890 50564
rect 2780 50244 2832 50250
rect 2780 50186 2832 50192
rect 2792 49978 2820 50186
rect 2780 49972 2832 49978
rect 2780 49914 2832 49920
rect 2582 49532 2890 49552
rect 2582 49530 2588 49532
rect 2644 49530 2668 49532
rect 2724 49530 2748 49532
rect 2804 49530 2828 49532
rect 2884 49530 2890 49532
rect 2644 49478 2646 49530
rect 2826 49478 2828 49530
rect 2582 49476 2588 49478
rect 2644 49476 2668 49478
rect 2724 49476 2748 49478
rect 2804 49476 2828 49478
rect 2884 49476 2890 49478
rect 2582 49456 2890 49476
rect 2688 49224 2740 49230
rect 2688 49166 2740 49172
rect 2700 48890 2728 49166
rect 2780 49088 2832 49094
rect 2780 49030 2832 49036
rect 2688 48884 2740 48890
rect 2688 48826 2740 48832
rect 2792 48793 2820 49030
rect 2778 48784 2834 48793
rect 2778 48719 2834 48728
rect 2582 48444 2890 48464
rect 2582 48442 2588 48444
rect 2644 48442 2668 48444
rect 2724 48442 2748 48444
rect 2804 48442 2828 48444
rect 2884 48442 2890 48444
rect 2644 48390 2646 48442
rect 2826 48390 2828 48442
rect 2582 48388 2588 48390
rect 2644 48388 2668 48390
rect 2724 48388 2748 48390
rect 2804 48388 2828 48390
rect 2884 48388 2890 48390
rect 2582 48368 2890 48388
rect 2688 48272 2740 48278
rect 2686 48240 2688 48249
rect 2740 48240 2742 48249
rect 2686 48175 2742 48184
rect 2976 47802 3004 51274
rect 3068 51074 3096 51342
rect 3344 51241 3372 54130
rect 3330 51232 3386 51241
rect 3330 51167 3386 51176
rect 3068 51046 3188 51074
rect 3056 50992 3108 50998
rect 3054 50960 3056 50969
rect 3108 50960 3110 50969
rect 3054 50895 3110 50904
rect 3056 50856 3108 50862
rect 3056 50798 3108 50804
rect 3068 50386 3096 50798
rect 3056 50380 3108 50386
rect 3056 50322 3108 50328
rect 3056 50244 3108 50250
rect 3056 50186 3108 50192
rect 2964 47796 3016 47802
rect 2964 47738 3016 47744
rect 2582 47356 2890 47376
rect 2582 47354 2588 47356
rect 2644 47354 2668 47356
rect 2724 47354 2748 47356
rect 2804 47354 2828 47356
rect 2884 47354 2890 47356
rect 2644 47302 2646 47354
rect 2826 47302 2828 47354
rect 2582 47300 2588 47302
rect 2644 47300 2668 47302
rect 2724 47300 2748 47302
rect 2804 47300 2828 47302
rect 2884 47300 2890 47302
rect 2582 47280 2890 47300
rect 2964 46912 3016 46918
rect 2964 46854 3016 46860
rect 2596 46708 2648 46714
rect 2596 46650 2648 46656
rect 2608 46578 2636 46650
rect 2976 46578 3004 46854
rect 3068 46753 3096 50186
rect 3160 48006 3188 51046
rect 3240 51060 3292 51066
rect 3240 51002 3292 51008
rect 3252 50946 3280 51002
rect 3436 50946 3464 61134
rect 3528 60602 3556 62070
rect 3620 60722 3648 66438
rect 3712 61674 3740 69702
rect 3792 68672 3844 68678
rect 3792 68614 3844 68620
rect 3804 67930 3832 68614
rect 3792 67924 3844 67930
rect 3792 67866 3844 67872
rect 3896 67658 3924 74802
rect 4620 74724 4672 74730
rect 4620 74666 4672 74672
rect 4213 74012 4521 74032
rect 4213 74010 4219 74012
rect 4275 74010 4299 74012
rect 4355 74010 4379 74012
rect 4435 74010 4459 74012
rect 4515 74010 4521 74012
rect 4275 73958 4277 74010
rect 4457 73958 4459 74010
rect 4213 73956 4219 73958
rect 4275 73956 4299 73958
rect 4355 73956 4379 73958
rect 4435 73956 4459 73958
rect 4515 73956 4521 73958
rect 4213 73936 4521 73956
rect 4213 72924 4521 72944
rect 4213 72922 4219 72924
rect 4275 72922 4299 72924
rect 4355 72922 4379 72924
rect 4435 72922 4459 72924
rect 4515 72922 4521 72924
rect 4275 72870 4277 72922
rect 4457 72870 4459 72922
rect 4213 72868 4219 72870
rect 4275 72868 4299 72870
rect 4355 72868 4379 72870
rect 4435 72868 4459 72870
rect 4515 72868 4521 72870
rect 4213 72848 4521 72868
rect 4213 71836 4521 71856
rect 4213 71834 4219 71836
rect 4275 71834 4299 71836
rect 4355 71834 4379 71836
rect 4435 71834 4459 71836
rect 4515 71834 4521 71836
rect 4275 71782 4277 71834
rect 4457 71782 4459 71834
rect 4213 71780 4219 71782
rect 4275 71780 4299 71782
rect 4355 71780 4379 71782
rect 4435 71780 4459 71782
rect 4515 71780 4521 71782
rect 4213 71760 4521 71780
rect 4068 70848 4120 70854
rect 4068 70790 4120 70796
rect 3976 69896 4028 69902
rect 3976 69838 4028 69844
rect 3988 69329 4016 69838
rect 3974 69320 4030 69329
rect 3974 69255 4030 69264
rect 3976 68808 4028 68814
rect 3976 68750 4028 68756
rect 3988 68513 4016 68750
rect 3974 68504 4030 68513
rect 3974 68439 4030 68448
rect 3884 67652 3936 67658
rect 3884 67594 3936 67600
rect 3792 64320 3844 64326
rect 3792 64262 3844 64268
rect 3700 61668 3752 61674
rect 3700 61610 3752 61616
rect 3608 60716 3660 60722
rect 3608 60658 3660 60664
rect 3528 60574 3740 60602
rect 3516 60512 3568 60518
rect 3516 60454 3568 60460
rect 3608 60512 3660 60518
rect 3608 60454 3660 60460
rect 3252 50918 3464 50946
rect 3330 50824 3386 50833
rect 3330 50759 3386 50768
rect 3240 50516 3292 50522
rect 3240 50458 3292 50464
rect 3252 50318 3280 50458
rect 3240 50312 3292 50318
rect 3240 50254 3292 50260
rect 3240 50176 3292 50182
rect 3240 50118 3292 50124
rect 3252 48142 3280 50118
rect 3240 48136 3292 48142
rect 3240 48078 3292 48084
rect 3148 48000 3200 48006
rect 3148 47942 3200 47948
rect 3148 47660 3200 47666
rect 3148 47602 3200 47608
rect 3054 46744 3110 46753
rect 3054 46679 3110 46688
rect 2596 46572 2648 46578
rect 2596 46514 2648 46520
rect 2964 46572 3016 46578
rect 3016 46532 3096 46560
rect 2964 46514 3016 46520
rect 2582 46268 2890 46288
rect 2582 46266 2588 46268
rect 2644 46266 2668 46268
rect 2724 46266 2748 46268
rect 2804 46266 2828 46268
rect 2884 46266 2890 46268
rect 2644 46214 2646 46266
rect 2826 46214 2828 46266
rect 2582 46212 2588 46214
rect 2644 46212 2668 46214
rect 2724 46212 2748 46214
rect 2804 46212 2828 46214
rect 2884 46212 2890 46214
rect 2582 46192 2890 46212
rect 2964 45824 3016 45830
rect 2962 45792 2964 45801
rect 3016 45792 3018 45801
rect 2962 45727 3018 45736
rect 2582 45180 2890 45200
rect 2582 45178 2588 45180
rect 2644 45178 2668 45180
rect 2724 45178 2748 45180
rect 2804 45178 2828 45180
rect 2884 45178 2890 45180
rect 2644 45126 2646 45178
rect 2826 45126 2828 45178
rect 2582 45124 2588 45126
rect 2644 45124 2668 45126
rect 2724 45124 2748 45126
rect 2804 45124 2828 45126
rect 2884 45124 2890 45126
rect 2582 45104 2890 45124
rect 2964 44872 3016 44878
rect 2964 44814 3016 44820
rect 2582 44092 2890 44112
rect 2582 44090 2588 44092
rect 2644 44090 2668 44092
rect 2724 44090 2748 44092
rect 2804 44090 2828 44092
rect 2884 44090 2890 44092
rect 2644 44038 2646 44090
rect 2826 44038 2828 44090
rect 2582 44036 2588 44038
rect 2644 44036 2668 44038
rect 2724 44036 2748 44038
rect 2804 44036 2828 44038
rect 2884 44036 2890 44038
rect 2582 44016 2890 44036
rect 2870 43344 2926 43353
rect 2870 43279 2926 43288
rect 2884 43246 2912 43279
rect 2872 43240 2924 43246
rect 2872 43182 2924 43188
rect 2582 43004 2890 43024
rect 2582 43002 2588 43004
rect 2644 43002 2668 43004
rect 2724 43002 2748 43004
rect 2804 43002 2828 43004
rect 2884 43002 2890 43004
rect 2644 42950 2646 43002
rect 2826 42950 2828 43002
rect 2582 42948 2588 42950
rect 2644 42948 2668 42950
rect 2724 42948 2748 42950
rect 2804 42948 2828 42950
rect 2884 42948 2890 42950
rect 2582 42928 2890 42948
rect 2582 41916 2890 41936
rect 2582 41914 2588 41916
rect 2644 41914 2668 41916
rect 2724 41914 2748 41916
rect 2804 41914 2828 41916
rect 2884 41914 2890 41916
rect 2644 41862 2646 41914
rect 2826 41862 2828 41914
rect 2582 41860 2588 41862
rect 2644 41860 2668 41862
rect 2724 41860 2748 41862
rect 2804 41860 2828 41862
rect 2884 41860 2890 41862
rect 2582 41840 2890 41860
rect 2516 41386 2636 41414
rect 2608 41018 2636 41386
rect 2332 39494 2452 39522
rect 2516 40990 2636 41018
rect 2228 39296 2280 39302
rect 2228 39238 2280 39244
rect 2240 38457 2268 39238
rect 2226 38448 2282 38457
rect 2226 38383 2282 38392
rect 2148 38270 2268 38298
rect 2240 38214 2268 38270
rect 2136 38208 2188 38214
rect 2136 38150 2188 38156
rect 2228 38208 2280 38214
rect 2228 38150 2280 38156
rect 2148 37398 2176 38150
rect 2332 37754 2360 39494
rect 2412 39432 2464 39438
rect 2412 39374 2464 39380
rect 2424 39030 2452 39374
rect 2412 39024 2464 39030
rect 2412 38966 2464 38972
rect 2412 38888 2464 38894
rect 2412 38830 2464 38836
rect 2424 38729 2452 38830
rect 2410 38720 2466 38729
rect 2410 38655 2466 38664
rect 2228 37732 2280 37738
rect 2332 37726 2452 37754
rect 2228 37674 2280 37680
rect 2136 37392 2188 37398
rect 2136 37334 2188 37340
rect 2136 37256 2188 37262
rect 2136 37198 2188 37204
rect 2044 32904 2096 32910
rect 2044 32846 2096 32852
rect 2148 32722 2176 37198
rect 2240 36786 2268 37674
rect 2318 37632 2374 37641
rect 2318 37567 2374 37576
rect 2332 37466 2360 37567
rect 2320 37460 2372 37466
rect 2320 37402 2372 37408
rect 2320 37324 2372 37330
rect 2320 37266 2372 37272
rect 2228 36780 2280 36786
rect 2228 36722 2280 36728
rect 2228 36576 2280 36582
rect 2228 36518 2280 36524
rect 2240 36281 2268 36518
rect 2226 36272 2282 36281
rect 2226 36207 2282 36216
rect 2332 35766 2360 37266
rect 2424 35873 2452 37726
rect 2410 35864 2466 35873
rect 2410 35799 2466 35808
rect 2320 35760 2372 35766
rect 2320 35702 2372 35708
rect 2228 34604 2280 34610
rect 2228 34546 2280 34552
rect 2240 34202 2268 34546
rect 2228 34196 2280 34202
rect 2228 34138 2280 34144
rect 2332 33946 2360 35702
rect 2412 35692 2464 35698
rect 2412 35634 2464 35640
rect 2424 35086 2452 35634
rect 2412 35080 2464 35086
rect 2412 35022 2464 35028
rect 2424 34610 2452 35022
rect 2412 34604 2464 34610
rect 2412 34546 2464 34552
rect 2240 33918 2360 33946
rect 2240 33538 2268 33918
rect 2320 33856 2372 33862
rect 2320 33798 2372 33804
rect 2332 33697 2360 33798
rect 2318 33688 2374 33697
rect 2318 33623 2374 33632
rect 2240 33510 2360 33538
rect 2424 33522 2452 34546
rect 2516 33522 2544 40990
rect 2582 40828 2890 40848
rect 2582 40826 2588 40828
rect 2644 40826 2668 40828
rect 2724 40826 2748 40828
rect 2804 40826 2828 40828
rect 2884 40826 2890 40828
rect 2644 40774 2646 40826
rect 2826 40774 2828 40826
rect 2582 40772 2588 40774
rect 2644 40772 2668 40774
rect 2724 40772 2748 40774
rect 2804 40772 2828 40774
rect 2884 40772 2890 40774
rect 2582 40752 2890 40772
rect 2780 40588 2832 40594
rect 2780 40530 2832 40536
rect 2792 40118 2820 40530
rect 2780 40112 2832 40118
rect 2780 40054 2832 40060
rect 2872 40044 2924 40050
rect 2872 39986 2924 39992
rect 2884 39914 2912 39986
rect 2872 39908 2924 39914
rect 2872 39850 2924 39856
rect 2582 39740 2890 39760
rect 2582 39738 2588 39740
rect 2644 39738 2668 39740
rect 2724 39738 2748 39740
rect 2804 39738 2828 39740
rect 2884 39738 2890 39740
rect 2644 39686 2646 39738
rect 2826 39686 2828 39738
rect 2582 39684 2588 39686
rect 2644 39684 2668 39686
rect 2724 39684 2748 39686
rect 2804 39684 2828 39686
rect 2884 39684 2890 39686
rect 2582 39664 2890 39684
rect 2976 39386 3004 44814
rect 3068 44402 3096 46532
rect 3056 44396 3108 44402
rect 3056 44338 3108 44344
rect 3056 43648 3108 43654
rect 3054 43616 3056 43625
rect 3108 43616 3110 43625
rect 3054 43551 3110 43560
rect 3054 43344 3110 43353
rect 3054 43279 3110 43288
rect 3068 40594 3096 43279
rect 3056 40588 3108 40594
rect 3056 40530 3108 40536
rect 3056 40384 3108 40390
rect 3056 40326 3108 40332
rect 3068 40225 3096 40326
rect 3054 40216 3110 40225
rect 3054 40151 3110 40160
rect 2976 39358 3096 39386
rect 2964 39296 3016 39302
rect 2964 39238 3016 39244
rect 2780 38956 2832 38962
rect 2780 38898 2832 38904
rect 2872 38956 2924 38962
rect 2872 38898 2924 38904
rect 2792 38826 2820 38898
rect 2780 38820 2832 38826
rect 2780 38762 2832 38768
rect 2884 38740 2912 38898
rect 2976 38865 3004 39238
rect 2962 38856 3018 38865
rect 2962 38791 3018 38800
rect 2884 38729 3004 38740
rect 2884 38720 3018 38729
rect 2884 38712 2962 38720
rect 2582 38652 2890 38672
rect 2962 38655 3018 38664
rect 2582 38650 2588 38652
rect 2644 38650 2668 38652
rect 2724 38650 2748 38652
rect 2804 38650 2828 38652
rect 2884 38650 2890 38652
rect 2644 38598 2646 38650
rect 2826 38598 2828 38650
rect 2582 38596 2588 38598
rect 2644 38596 2668 38598
rect 2724 38596 2748 38598
rect 2804 38596 2828 38598
rect 2884 38596 2890 38598
rect 2582 38576 2890 38596
rect 2780 38344 2832 38350
rect 2780 38286 2832 38292
rect 2792 37874 2820 38286
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2582 37564 2890 37584
rect 2582 37562 2588 37564
rect 2644 37562 2668 37564
rect 2724 37562 2748 37564
rect 2804 37562 2828 37564
rect 2884 37562 2890 37564
rect 2644 37510 2646 37562
rect 2826 37510 2828 37562
rect 2582 37508 2588 37510
rect 2644 37508 2668 37510
rect 2724 37508 2748 37510
rect 2804 37508 2828 37510
rect 2884 37508 2890 37510
rect 2582 37488 2890 37508
rect 2976 37233 3004 38655
rect 2962 37224 3018 37233
rect 2962 37159 3018 37168
rect 2780 37120 2832 37126
rect 3068 37074 3096 39358
rect 2780 37062 2832 37068
rect 2792 36786 2820 37062
rect 2976 37046 3096 37074
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2582 36476 2890 36496
rect 2582 36474 2588 36476
rect 2644 36474 2668 36476
rect 2724 36474 2748 36476
rect 2804 36474 2828 36476
rect 2884 36474 2890 36476
rect 2644 36422 2646 36474
rect 2826 36422 2828 36474
rect 2582 36420 2588 36422
rect 2644 36420 2668 36422
rect 2724 36420 2748 36422
rect 2804 36420 2828 36422
rect 2884 36420 2890 36422
rect 2582 36400 2890 36420
rect 2582 35388 2890 35408
rect 2582 35386 2588 35388
rect 2644 35386 2668 35388
rect 2724 35386 2748 35388
rect 2804 35386 2828 35388
rect 2884 35386 2890 35388
rect 2644 35334 2646 35386
rect 2826 35334 2828 35386
rect 2582 35332 2588 35334
rect 2644 35332 2668 35334
rect 2724 35332 2748 35334
rect 2804 35332 2828 35334
rect 2884 35332 2890 35334
rect 2582 35312 2890 35332
rect 2582 34300 2890 34320
rect 2582 34298 2588 34300
rect 2644 34298 2668 34300
rect 2724 34298 2748 34300
rect 2804 34298 2828 34300
rect 2884 34298 2890 34300
rect 2644 34246 2646 34298
rect 2826 34246 2828 34298
rect 2582 34244 2588 34246
rect 2644 34244 2668 34246
rect 2724 34244 2748 34246
rect 2804 34244 2828 34246
rect 2884 34244 2890 34246
rect 2582 34224 2890 34244
rect 2228 33448 2280 33454
rect 2228 33390 2280 33396
rect 2056 32694 2176 32722
rect 1952 32496 2004 32502
rect 1952 32438 2004 32444
rect 1860 30320 1912 30326
rect 1860 30262 1912 30268
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1872 29458 1900 30126
rect 1688 29430 1900 29458
rect 1584 26444 1636 26450
rect 1584 26386 1636 26392
rect 1492 26376 1544 26382
rect 1492 26318 1544 26324
rect 1398 25936 1454 25945
rect 1398 25871 1454 25880
rect 1504 25537 1532 26318
rect 1584 26240 1636 26246
rect 1584 26182 1636 26188
rect 1490 25528 1546 25537
rect 1490 25463 1546 25472
rect 1492 24812 1544 24818
rect 1492 24754 1544 24760
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 22953 1440 24142
rect 1504 23361 1532 24754
rect 1596 24206 1624 26182
rect 1584 24200 1636 24206
rect 1584 24142 1636 24148
rect 1584 23520 1636 23526
rect 1584 23462 1636 23468
rect 1490 23352 1546 23361
rect 1490 23287 1546 23296
rect 1596 23118 1624 23462
rect 1584 23112 1636 23118
rect 1584 23054 1636 23060
rect 1398 22944 1454 22953
rect 1398 22879 1454 22888
rect 1688 20602 1716 29430
rect 1766 29200 1822 29209
rect 1766 29135 1822 29144
rect 1780 21690 1808 29135
rect 1964 27878 1992 32438
rect 2056 30122 2084 32694
rect 2136 32428 2188 32434
rect 2136 32370 2188 32376
rect 2148 30394 2176 32370
rect 2240 31793 2268 33390
rect 2332 32978 2360 33510
rect 2412 33516 2464 33522
rect 2412 33458 2464 33464
rect 2504 33516 2556 33522
rect 2504 33458 2556 33464
rect 2582 33212 2890 33232
rect 2582 33210 2588 33212
rect 2644 33210 2668 33212
rect 2724 33210 2748 33212
rect 2804 33210 2828 33212
rect 2884 33210 2890 33212
rect 2644 33158 2646 33210
rect 2826 33158 2828 33210
rect 2582 33156 2588 33158
rect 2644 33156 2668 33158
rect 2724 33156 2748 33158
rect 2804 33156 2828 33158
rect 2884 33156 2890 33158
rect 2582 33136 2890 33156
rect 2976 33114 3004 37046
rect 3054 36680 3110 36689
rect 3054 36615 3056 36624
rect 3108 36615 3110 36624
rect 3056 36586 3108 36592
rect 3054 34504 3110 34513
rect 3054 34439 3110 34448
rect 3068 34134 3096 34439
rect 3056 34128 3108 34134
rect 3056 34070 3108 34076
rect 2964 33108 3016 33114
rect 2964 33050 3016 33056
rect 2320 32972 2372 32978
rect 2320 32914 2372 32920
rect 2504 32972 2556 32978
rect 2504 32914 2556 32920
rect 2318 32872 2374 32881
rect 2318 32807 2374 32816
rect 2332 32774 2360 32807
rect 2320 32768 2372 32774
rect 2320 32710 2372 32716
rect 2318 32600 2374 32609
rect 2516 32570 2544 32914
rect 2318 32535 2374 32544
rect 2504 32564 2556 32570
rect 2332 32230 2360 32535
rect 2504 32506 2556 32512
rect 2502 32464 2558 32473
rect 2502 32399 2558 32408
rect 2320 32224 2372 32230
rect 2320 32166 2372 32172
rect 2320 31884 2372 31890
rect 2320 31826 2372 31832
rect 2226 31784 2282 31793
rect 2226 31719 2282 31728
rect 2226 31648 2282 31657
rect 2226 31583 2282 31592
rect 2136 30388 2188 30394
rect 2136 30330 2188 30336
rect 2136 30252 2188 30258
rect 2136 30194 2188 30200
rect 2044 30116 2096 30122
rect 2044 30058 2096 30064
rect 2148 29345 2176 30194
rect 2134 29336 2190 29345
rect 2044 29300 2096 29306
rect 2134 29271 2190 29280
rect 2044 29242 2096 29248
rect 1952 27872 2004 27878
rect 1952 27814 2004 27820
rect 1860 27328 1912 27334
rect 1860 27270 1912 27276
rect 1872 25906 1900 27270
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 1964 26586 1992 26930
rect 1952 26580 2004 26586
rect 1952 26522 2004 26528
rect 1952 26444 2004 26450
rect 1952 26386 2004 26392
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1860 25764 1912 25770
rect 1860 25706 1912 25712
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1768 21480 1820 21486
rect 1768 21422 1820 21428
rect 1780 20806 1808 21422
rect 1768 20800 1820 20806
rect 1768 20742 1820 20748
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 17785 1440 19314
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 1596 17678 1624 19110
rect 1872 18426 1900 25706
rect 1964 21146 1992 26386
rect 2056 25786 2084 29242
rect 2136 27464 2188 27470
rect 2136 27406 2188 27412
rect 2148 26382 2176 27406
rect 2240 27010 2268 31583
rect 2332 30954 2360 31826
rect 2412 31680 2464 31686
rect 2412 31622 2464 31628
rect 2424 31521 2452 31622
rect 2410 31512 2466 31521
rect 2410 31447 2466 31456
rect 2412 31136 2464 31142
rect 2410 31104 2412 31113
rect 2464 31104 2466 31113
rect 2410 31039 2466 31048
rect 2332 30926 2452 30954
rect 2320 30728 2372 30734
rect 2320 30670 2372 30676
rect 2332 30297 2360 30670
rect 2318 30288 2374 30297
rect 2318 30223 2374 30232
rect 2424 29306 2452 30926
rect 2412 29300 2464 29306
rect 2412 29242 2464 29248
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 2424 29050 2452 29106
rect 2332 29022 2452 29050
rect 2332 28082 2360 29022
rect 2516 28994 2544 32399
rect 2582 32124 2890 32144
rect 2582 32122 2588 32124
rect 2644 32122 2668 32124
rect 2724 32122 2748 32124
rect 2804 32122 2828 32124
rect 2884 32122 2890 32124
rect 2644 32070 2646 32122
rect 2826 32070 2828 32122
rect 2582 32068 2588 32070
rect 2644 32068 2668 32070
rect 2724 32068 2748 32070
rect 2804 32068 2828 32070
rect 2884 32068 2890 32070
rect 2582 32048 2890 32068
rect 3056 31272 3108 31278
rect 3056 31214 3108 31220
rect 2582 31036 2890 31056
rect 2582 31034 2588 31036
rect 2644 31034 2668 31036
rect 2724 31034 2748 31036
rect 2804 31034 2828 31036
rect 2884 31034 2890 31036
rect 2644 30982 2646 31034
rect 2826 30982 2828 31034
rect 2582 30980 2588 30982
rect 2644 30980 2668 30982
rect 2724 30980 2748 30982
rect 2804 30980 2828 30982
rect 2884 30980 2890 30982
rect 2582 30960 2890 30980
rect 2964 30252 3016 30258
rect 2964 30194 3016 30200
rect 2582 29948 2890 29968
rect 2582 29946 2588 29948
rect 2644 29946 2668 29948
rect 2724 29946 2748 29948
rect 2804 29946 2828 29948
rect 2884 29946 2890 29948
rect 2644 29894 2646 29946
rect 2826 29894 2828 29946
rect 2582 29892 2588 29894
rect 2644 29892 2668 29894
rect 2724 29892 2748 29894
rect 2804 29892 2828 29894
rect 2884 29892 2890 29894
rect 2582 29872 2890 29892
rect 2976 29753 3004 30194
rect 3068 29850 3096 31214
rect 3056 29844 3108 29850
rect 3056 29786 3108 29792
rect 2962 29744 3018 29753
rect 2962 29679 3018 29688
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 3056 29640 3108 29646
rect 3056 29582 3108 29588
rect 2780 29232 2832 29238
rect 2780 29174 2832 29180
rect 2792 29017 2820 29174
rect 2424 28966 2544 28994
rect 2778 29008 2834 29017
rect 2424 28200 2452 28966
rect 2976 28966 3004 29582
rect 3068 28966 3096 29582
rect 2778 28943 2834 28952
rect 2964 28960 3016 28966
rect 2964 28902 3016 28908
rect 3056 28960 3108 28966
rect 3056 28902 3108 28908
rect 2582 28860 2890 28880
rect 2582 28858 2588 28860
rect 2644 28858 2668 28860
rect 2724 28858 2748 28860
rect 2804 28858 2828 28860
rect 2884 28858 2890 28860
rect 2644 28806 2646 28858
rect 2826 28806 2828 28858
rect 2582 28804 2588 28806
rect 2644 28804 2668 28806
rect 2724 28804 2748 28806
rect 2804 28804 2828 28806
rect 2884 28804 2890 28806
rect 2582 28784 2890 28804
rect 2780 28552 2832 28558
rect 2780 28494 2832 28500
rect 2688 28416 2740 28422
rect 2688 28358 2740 28364
rect 2424 28172 2544 28200
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2332 27470 2360 28018
rect 2424 27674 2452 28018
rect 2412 27668 2464 27674
rect 2412 27610 2464 27616
rect 2320 27464 2372 27470
rect 2320 27406 2372 27412
rect 2332 27130 2360 27406
rect 2320 27124 2372 27130
rect 2320 27066 2372 27072
rect 2240 26982 2360 27010
rect 2228 26920 2280 26926
rect 2228 26862 2280 26868
rect 2136 26376 2188 26382
rect 2136 26318 2188 26324
rect 2148 25945 2176 26318
rect 2134 25936 2190 25945
rect 2134 25871 2190 25880
rect 2056 25758 2176 25786
rect 2044 25696 2096 25702
rect 2044 25638 2096 25644
rect 2056 25294 2084 25638
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 2148 24154 2176 25758
rect 2056 24126 2176 24154
rect 1952 21140 2004 21146
rect 1952 21082 2004 21088
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1964 18850 1992 20742
rect 2056 18970 2084 24126
rect 2136 24064 2188 24070
rect 2136 24006 2188 24012
rect 2148 23118 2176 24006
rect 2136 23112 2188 23118
rect 2136 23054 2188 23060
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 1964 18822 2084 18850
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1860 18420 1912 18426
rect 1860 18362 1912 18368
rect 1964 18290 1992 18566
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1412 14958 1440 16390
rect 1492 16108 1544 16114
rect 1492 16050 1544 16056
rect 1504 15162 1532 16050
rect 1596 15502 1624 16934
rect 1780 16114 1808 16934
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15706 1716 15982
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1584 15496 1636 15502
rect 1584 15438 1636 15444
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 12345 1440 13262
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1228 11750 1348 11778
rect 1228 5302 1256 11750
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 10985 1348 11630
rect 1412 11393 1440 12174
rect 1504 11801 1532 12718
rect 1490 11792 1546 11801
rect 1490 11727 1546 11736
rect 1398 11384 1454 11393
rect 1398 11319 1454 11328
rect 1584 11280 1636 11286
rect 1584 11222 1636 11228
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1306 10976 1362 10985
rect 1306 10911 1362 10920
rect 1308 10600 1360 10606
rect 1308 10542 1360 10548
rect 1320 10033 1348 10542
rect 1412 10441 1440 11086
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1400 10056 1452 10062
rect 1306 10024 1362 10033
rect 1400 9998 1452 10004
rect 1306 9959 1362 9968
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9217 1440 9454
rect 1398 9208 1454 9217
rect 1596 9178 1624 11222
rect 1780 10674 1808 15438
rect 1872 15201 1900 16050
rect 1858 15192 1914 15201
rect 1858 15127 1914 15136
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1872 14618 1900 14962
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 13025 1900 13874
rect 1964 13394 1992 17478
rect 2056 16250 2084 18822
rect 2148 18222 2176 21626
rect 2240 19514 2268 26862
rect 2332 26330 2360 26982
rect 2424 26518 2452 27610
rect 2412 26512 2464 26518
rect 2412 26454 2464 26460
rect 2332 26302 2452 26330
rect 2320 26240 2372 26246
rect 2320 26182 2372 26188
rect 2332 25294 2360 26182
rect 2320 25288 2372 25294
rect 2320 25230 2372 25236
rect 2320 24948 2372 24954
rect 2320 24890 2372 24896
rect 2332 21690 2360 24890
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2332 21146 2360 21490
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2320 20460 2372 20466
rect 2320 20402 2372 20408
rect 2228 19508 2280 19514
rect 2332 19496 2360 20402
rect 2424 20058 2452 26302
rect 2516 24154 2544 28172
rect 2700 28150 2728 28358
rect 2792 28218 2820 28494
rect 2780 28212 2832 28218
rect 2780 28154 2832 28160
rect 2688 28144 2740 28150
rect 2688 28086 2740 28092
rect 3056 28076 3108 28082
rect 3056 28018 3108 28024
rect 2582 27772 2890 27792
rect 2582 27770 2588 27772
rect 2644 27770 2668 27772
rect 2724 27770 2748 27772
rect 2804 27770 2828 27772
rect 2884 27770 2890 27772
rect 2644 27718 2646 27770
rect 2826 27718 2828 27770
rect 2582 27716 2588 27718
rect 2644 27716 2668 27718
rect 2724 27716 2748 27718
rect 2804 27716 2828 27718
rect 2884 27716 2890 27718
rect 2582 27696 2890 27716
rect 2778 27568 2834 27577
rect 2778 27503 2834 27512
rect 2872 27532 2924 27538
rect 2596 27464 2648 27470
rect 2596 27406 2648 27412
rect 2608 26994 2636 27406
rect 2792 27402 2820 27503
rect 2872 27474 2924 27480
rect 2884 27441 2912 27474
rect 2870 27432 2926 27441
rect 2780 27396 2832 27402
rect 2870 27367 2926 27376
rect 2780 27338 2832 27344
rect 2872 27328 2924 27334
rect 2872 27270 2924 27276
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2884 26858 2912 27270
rect 3068 26994 3096 28018
rect 3056 26988 3108 26994
rect 3056 26930 3108 26936
rect 2872 26852 2924 26858
rect 2872 26794 2924 26800
rect 2582 26684 2890 26704
rect 2582 26682 2588 26684
rect 2644 26682 2668 26684
rect 2724 26682 2748 26684
rect 2804 26682 2828 26684
rect 2884 26682 2890 26684
rect 2644 26630 2646 26682
rect 2826 26630 2828 26682
rect 2582 26628 2588 26630
rect 2644 26628 2668 26630
rect 2724 26628 2748 26630
rect 2804 26628 2828 26630
rect 2884 26628 2890 26630
rect 2582 26608 2890 26628
rect 2596 26512 2648 26518
rect 2596 26454 2648 26460
rect 2608 25838 2636 26454
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2596 25832 2648 25838
rect 2596 25774 2648 25780
rect 2582 25596 2890 25616
rect 2582 25594 2588 25596
rect 2644 25594 2668 25596
rect 2724 25594 2748 25596
rect 2804 25594 2828 25596
rect 2884 25594 2890 25596
rect 2644 25542 2646 25594
rect 2826 25542 2828 25594
rect 2582 25540 2588 25542
rect 2644 25540 2668 25542
rect 2724 25540 2748 25542
rect 2804 25540 2828 25542
rect 2884 25540 2890 25542
rect 2582 25520 2890 25540
rect 2594 25392 2650 25401
rect 2594 25327 2650 25336
rect 2608 24954 2636 25327
rect 2872 25152 2924 25158
rect 2976 25129 3004 25842
rect 2872 25094 2924 25100
rect 2962 25120 3018 25129
rect 2596 24948 2648 24954
rect 2596 24890 2648 24896
rect 2884 24818 2912 25094
rect 2962 25055 3018 25064
rect 2872 24812 2924 24818
rect 2872 24754 2924 24760
rect 2964 24676 3016 24682
rect 2964 24618 3016 24624
rect 2582 24508 2890 24528
rect 2582 24506 2588 24508
rect 2644 24506 2668 24508
rect 2724 24506 2748 24508
rect 2804 24506 2828 24508
rect 2884 24506 2890 24508
rect 2644 24454 2646 24506
rect 2826 24454 2828 24506
rect 2582 24452 2588 24454
rect 2644 24452 2668 24454
rect 2724 24452 2748 24454
rect 2804 24452 2828 24454
rect 2884 24452 2890 24454
rect 2582 24432 2890 24452
rect 2516 24126 2636 24154
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2516 23730 2544 24006
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2608 23508 2636 24126
rect 2516 23480 2636 23508
rect 2516 23322 2544 23480
rect 2582 23420 2890 23440
rect 2582 23418 2588 23420
rect 2644 23418 2668 23420
rect 2724 23418 2748 23420
rect 2804 23418 2828 23420
rect 2884 23418 2890 23420
rect 2644 23366 2646 23418
rect 2826 23366 2828 23418
rect 2582 23364 2588 23366
rect 2644 23364 2668 23366
rect 2724 23364 2748 23366
rect 2804 23364 2828 23366
rect 2884 23364 2890 23366
rect 2582 23344 2890 23364
rect 2504 23316 2556 23322
rect 2504 23258 2556 23264
rect 2976 23118 3004 24618
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2582 22332 2890 22352
rect 2582 22330 2588 22332
rect 2644 22330 2668 22332
rect 2724 22330 2748 22332
rect 2804 22330 2828 22332
rect 2884 22330 2890 22332
rect 2644 22278 2646 22330
rect 2826 22278 2828 22330
rect 2582 22276 2588 22278
rect 2644 22276 2668 22278
rect 2724 22276 2748 22278
rect 2804 22276 2828 22278
rect 2884 22276 2890 22278
rect 2582 22256 2890 22276
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2884 21457 2912 21966
rect 2870 21448 2926 21457
rect 2504 21412 2556 21418
rect 2870 21383 2926 21392
rect 2504 21354 2556 21360
rect 2516 20874 2544 21354
rect 2582 21244 2890 21264
rect 2582 21242 2588 21244
rect 2644 21242 2668 21244
rect 2724 21242 2748 21244
rect 2804 21242 2828 21244
rect 2884 21242 2890 21244
rect 2644 21190 2646 21242
rect 2826 21190 2828 21242
rect 2582 21188 2588 21190
rect 2644 21188 2668 21190
rect 2724 21188 2748 21190
rect 2804 21188 2828 21190
rect 2884 21188 2890 21190
rect 2582 21168 2890 21188
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2412 19508 2464 19514
rect 2332 19468 2412 19496
rect 2228 19450 2280 19456
rect 2412 19450 2464 19456
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15570 2084 15846
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2148 15450 2176 17614
rect 2240 17338 2268 18226
rect 2332 17678 2360 18634
rect 2424 18426 2452 19314
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2240 16561 2268 17138
rect 2226 16552 2282 16561
rect 2226 16487 2282 16496
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 15570 2360 16458
rect 2516 16454 2544 20810
rect 2792 20466 2820 21014
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2582 20156 2890 20176
rect 2582 20154 2588 20156
rect 2644 20154 2668 20156
rect 2724 20154 2748 20156
rect 2804 20154 2828 20156
rect 2884 20154 2890 20156
rect 2644 20102 2646 20154
rect 2826 20102 2828 20154
rect 2582 20100 2588 20102
rect 2644 20100 2668 20102
rect 2724 20100 2748 20102
rect 2804 20100 2828 20102
rect 2884 20100 2890 20102
rect 2582 20080 2890 20100
rect 2582 19068 2890 19088
rect 2582 19066 2588 19068
rect 2644 19066 2668 19068
rect 2724 19066 2748 19068
rect 2804 19066 2828 19068
rect 2884 19066 2890 19068
rect 2644 19014 2646 19066
rect 2826 19014 2828 19066
rect 2582 19012 2588 19014
rect 2644 19012 2668 19014
rect 2724 19012 2748 19014
rect 2804 19012 2828 19014
rect 2884 19012 2890 19014
rect 2582 18992 2890 19012
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2792 18193 2820 18702
rect 2778 18184 2834 18193
rect 2778 18119 2834 18128
rect 2582 17980 2890 18000
rect 2582 17978 2588 17980
rect 2644 17978 2668 17980
rect 2724 17978 2748 17980
rect 2804 17978 2828 17980
rect 2884 17978 2890 17980
rect 2644 17926 2646 17978
rect 2826 17926 2828 17978
rect 2582 17924 2588 17926
rect 2644 17924 2668 17926
rect 2724 17924 2748 17926
rect 2804 17924 2828 17926
rect 2884 17924 2890 17926
rect 2582 17904 2890 17924
rect 2976 17746 3004 20742
rect 3068 20602 3096 26930
rect 3160 24290 3188 47602
rect 3252 46578 3280 48078
rect 3240 46572 3292 46578
rect 3240 46514 3292 46520
rect 3240 46436 3292 46442
rect 3240 46378 3292 46384
rect 3252 44742 3280 46378
rect 3240 44736 3292 44742
rect 3240 44678 3292 44684
rect 3344 44538 3372 50759
rect 3424 50244 3476 50250
rect 3424 50186 3476 50192
rect 3436 45665 3464 50186
rect 3422 45656 3478 45665
rect 3422 45591 3478 45600
rect 3424 45416 3476 45422
rect 3424 45358 3476 45364
rect 3332 44532 3384 44538
rect 3332 44474 3384 44480
rect 3240 44396 3292 44402
rect 3240 44338 3292 44344
rect 3252 41614 3280 44338
rect 3332 44328 3384 44334
rect 3332 44270 3384 44276
rect 3344 43314 3372 44270
rect 3436 43790 3464 45358
rect 3424 43784 3476 43790
rect 3424 43726 3476 43732
rect 3332 43308 3384 43314
rect 3332 43250 3384 43256
rect 3332 42900 3384 42906
rect 3332 42842 3384 42848
rect 3344 42106 3372 42842
rect 3436 42294 3464 43726
rect 3424 42288 3476 42294
rect 3424 42230 3476 42236
rect 3344 42078 3464 42106
rect 3240 41608 3292 41614
rect 3240 41550 3292 41556
rect 3332 40656 3384 40662
rect 3332 40598 3384 40604
rect 3240 40112 3292 40118
rect 3240 40054 3292 40060
rect 3252 38554 3280 40054
rect 3240 38548 3292 38554
rect 3240 38490 3292 38496
rect 3240 38412 3292 38418
rect 3240 38354 3292 38360
rect 3252 34610 3280 38354
rect 3240 34604 3292 34610
rect 3240 34546 3292 34552
rect 3240 34400 3292 34406
rect 3240 34342 3292 34348
rect 3252 34105 3280 34342
rect 3238 34096 3294 34105
rect 3238 34031 3294 34040
rect 3344 33998 3372 40598
rect 3436 37262 3464 42078
rect 3528 40662 3556 60454
rect 3620 56506 3648 60454
rect 3712 57633 3740 60574
rect 3698 57624 3754 57633
rect 3698 57559 3754 57568
rect 3700 57316 3752 57322
rect 3700 57258 3752 57264
rect 3608 56500 3660 56506
rect 3608 56442 3660 56448
rect 3608 56296 3660 56302
rect 3608 56238 3660 56244
rect 3620 44538 3648 56238
rect 3712 51542 3740 57258
rect 3804 51610 3832 64262
rect 3882 63880 3938 63889
rect 3882 63815 3884 63824
rect 3936 63815 3938 63824
rect 3884 63786 3936 63792
rect 4080 63481 4108 70790
rect 4213 70748 4521 70768
rect 4213 70746 4219 70748
rect 4275 70746 4299 70748
rect 4355 70746 4379 70748
rect 4435 70746 4459 70748
rect 4515 70746 4521 70748
rect 4275 70694 4277 70746
rect 4457 70694 4459 70746
rect 4213 70692 4219 70694
rect 4275 70692 4299 70694
rect 4355 70692 4379 70694
rect 4435 70692 4459 70694
rect 4515 70692 4521 70694
rect 4213 70672 4521 70692
rect 4213 69660 4521 69680
rect 4213 69658 4219 69660
rect 4275 69658 4299 69660
rect 4355 69658 4379 69660
rect 4435 69658 4459 69660
rect 4515 69658 4521 69660
rect 4275 69606 4277 69658
rect 4457 69606 4459 69658
rect 4213 69604 4219 69606
rect 4275 69604 4299 69606
rect 4355 69604 4379 69606
rect 4435 69604 4459 69606
rect 4515 69604 4521 69606
rect 4213 69584 4521 69604
rect 4160 69420 4212 69426
rect 4160 69362 4212 69368
rect 4172 68921 4200 69362
rect 4158 68912 4214 68921
rect 4158 68847 4214 68856
rect 4213 68572 4521 68592
rect 4213 68570 4219 68572
rect 4275 68570 4299 68572
rect 4355 68570 4379 68572
rect 4435 68570 4459 68572
rect 4515 68570 4521 68572
rect 4275 68518 4277 68570
rect 4457 68518 4459 68570
rect 4213 68516 4219 68518
rect 4275 68516 4299 68518
rect 4355 68516 4379 68518
rect 4435 68516 4459 68518
rect 4515 68516 4521 68518
rect 4213 68496 4521 68516
rect 4213 67484 4521 67504
rect 4213 67482 4219 67484
rect 4275 67482 4299 67484
rect 4355 67482 4379 67484
rect 4435 67482 4459 67484
rect 4515 67482 4521 67484
rect 4275 67430 4277 67482
rect 4457 67430 4459 67482
rect 4213 67428 4219 67430
rect 4275 67428 4299 67430
rect 4355 67428 4379 67430
rect 4435 67428 4459 67430
rect 4515 67428 4521 67430
rect 4213 67408 4521 67428
rect 4213 66396 4521 66416
rect 4213 66394 4219 66396
rect 4275 66394 4299 66396
rect 4355 66394 4379 66396
rect 4435 66394 4459 66396
rect 4515 66394 4521 66396
rect 4275 66342 4277 66394
rect 4457 66342 4459 66394
rect 4213 66340 4219 66342
rect 4275 66340 4299 66342
rect 4355 66340 4379 66342
rect 4435 66340 4459 66342
rect 4515 66340 4521 66342
rect 4213 66320 4521 66340
rect 4213 65308 4521 65328
rect 4213 65306 4219 65308
rect 4275 65306 4299 65308
rect 4355 65306 4379 65308
rect 4435 65306 4459 65308
rect 4515 65306 4521 65308
rect 4275 65254 4277 65306
rect 4457 65254 4459 65306
rect 4213 65252 4219 65254
rect 4275 65252 4299 65254
rect 4355 65252 4379 65254
rect 4435 65252 4459 65254
rect 4515 65252 4521 65254
rect 4213 65232 4521 65252
rect 4213 64220 4521 64240
rect 4213 64218 4219 64220
rect 4275 64218 4299 64220
rect 4355 64218 4379 64220
rect 4435 64218 4459 64220
rect 4515 64218 4521 64220
rect 4275 64166 4277 64218
rect 4457 64166 4459 64218
rect 4213 64164 4219 64166
rect 4275 64164 4299 64166
rect 4355 64164 4379 64166
rect 4435 64164 4459 64166
rect 4515 64164 4521 64166
rect 4213 64144 4521 64164
rect 4066 63472 4122 63481
rect 4066 63407 4122 63416
rect 3884 63300 3936 63306
rect 3884 63242 3936 63248
rect 4068 63300 4120 63306
rect 4068 63242 4120 63248
rect 3896 62286 3924 63242
rect 3976 63232 4028 63238
rect 4080 63209 4108 63242
rect 3976 63174 4028 63180
rect 4066 63200 4122 63209
rect 3988 62937 4016 63174
rect 4066 63135 4122 63144
rect 4213 63132 4521 63152
rect 4213 63130 4219 63132
rect 4275 63130 4299 63132
rect 4355 63130 4379 63132
rect 4435 63130 4459 63132
rect 4515 63130 4521 63132
rect 4275 63078 4277 63130
rect 4457 63078 4459 63130
rect 4213 63076 4219 63078
rect 4275 63076 4299 63078
rect 4355 63076 4379 63078
rect 4435 63076 4459 63078
rect 4515 63076 4521 63078
rect 4213 63056 4521 63076
rect 3974 62928 4030 62937
rect 3974 62863 4030 62872
rect 3884 62280 3936 62286
rect 3884 62222 3936 62228
rect 3896 60761 3924 62222
rect 4213 62044 4521 62064
rect 4213 62042 4219 62044
rect 4275 62042 4299 62044
rect 4355 62042 4379 62044
rect 4435 62042 4459 62044
rect 4515 62042 4521 62044
rect 4275 61990 4277 62042
rect 4457 61990 4459 62042
rect 4213 61988 4219 61990
rect 4275 61988 4299 61990
rect 4355 61988 4379 61990
rect 4435 61988 4459 61990
rect 4515 61988 4521 61990
rect 4213 61968 4521 61988
rect 4068 61940 4120 61946
rect 4068 61882 4120 61888
rect 3974 61160 4030 61169
rect 3974 61095 4030 61104
rect 3988 61062 4016 61095
rect 3976 61056 4028 61062
rect 3976 60998 4028 61004
rect 3882 60752 3938 60761
rect 3882 60687 3938 60696
rect 3976 60308 4028 60314
rect 3976 60250 4028 60256
rect 3988 56302 4016 60250
rect 3976 56296 4028 56302
rect 3976 56238 4028 56244
rect 3976 55616 4028 55622
rect 3974 55584 3976 55593
rect 4028 55584 4030 55593
rect 3974 55519 4030 55528
rect 3976 55344 4028 55350
rect 3976 55286 4028 55292
rect 3792 51604 3844 51610
rect 3792 51546 3844 51552
rect 3700 51536 3752 51542
rect 3700 51478 3752 51484
rect 3698 51096 3754 51105
rect 3698 51031 3700 51040
rect 3752 51031 3754 51040
rect 3700 51002 3752 51008
rect 3700 50924 3752 50930
rect 3700 50866 3752 50872
rect 3712 50182 3740 50866
rect 3790 50552 3846 50561
rect 3790 50487 3846 50496
rect 3700 50176 3752 50182
rect 3700 50118 3752 50124
rect 3700 49836 3752 49842
rect 3700 49778 3752 49784
rect 3712 49162 3740 49778
rect 3700 49156 3752 49162
rect 3700 49098 3752 49104
rect 3712 48754 3740 49098
rect 3700 48748 3752 48754
rect 3700 48690 3752 48696
rect 3712 45422 3740 48690
rect 3804 47258 3832 50487
rect 3884 50312 3936 50318
rect 3884 50254 3936 50260
rect 3896 49842 3924 50254
rect 3884 49836 3936 49842
rect 3884 49778 3936 49784
rect 3882 49600 3938 49609
rect 3882 49535 3938 49544
rect 3896 49298 3924 49535
rect 3884 49292 3936 49298
rect 3884 49234 3936 49240
rect 3882 49192 3938 49201
rect 3882 49127 3938 49136
rect 3792 47252 3844 47258
rect 3792 47194 3844 47200
rect 3896 47138 3924 49127
rect 3804 47110 3924 47138
rect 3700 45416 3752 45422
rect 3700 45358 3752 45364
rect 3712 44878 3740 45358
rect 3804 44985 3832 47110
rect 3884 46572 3936 46578
rect 3884 46514 3936 46520
rect 3790 44976 3846 44985
rect 3790 44911 3846 44920
rect 3700 44872 3752 44878
rect 3700 44814 3752 44820
rect 3792 44872 3844 44878
rect 3792 44814 3844 44820
rect 3700 44736 3752 44742
rect 3700 44678 3752 44684
rect 3608 44532 3660 44538
rect 3608 44474 3660 44480
rect 3606 44432 3662 44441
rect 3606 44367 3662 44376
rect 3620 43858 3648 44367
rect 3608 43852 3660 43858
rect 3608 43794 3660 43800
rect 3608 42288 3660 42294
rect 3608 42230 3660 42236
rect 3516 40656 3568 40662
rect 3516 40598 3568 40604
rect 3516 40520 3568 40526
rect 3516 40462 3568 40468
rect 3528 40050 3556 40462
rect 3516 40044 3568 40050
rect 3516 39986 3568 39992
rect 3514 39944 3570 39953
rect 3514 39879 3570 39888
rect 3528 38486 3556 39879
rect 3620 38826 3648 42230
rect 3712 41478 3740 44678
rect 3804 44402 3832 44814
rect 3792 44396 3844 44402
rect 3792 44338 3844 44344
rect 3896 44266 3924 46514
rect 3884 44260 3936 44266
rect 3884 44202 3936 44208
rect 3988 42786 4016 55286
rect 3804 42758 4016 42786
rect 3700 41472 3752 41478
rect 3700 41414 3752 41420
rect 3804 40730 3832 42758
rect 3976 42084 4028 42090
rect 3976 42026 4028 42032
rect 3792 40724 3844 40730
rect 3792 40666 3844 40672
rect 3700 40452 3752 40458
rect 3700 40394 3752 40400
rect 3712 39030 3740 40394
rect 3988 40118 4016 42026
rect 3976 40112 4028 40118
rect 4080 40089 4108 61882
rect 4213 60956 4521 60976
rect 4213 60954 4219 60956
rect 4275 60954 4299 60956
rect 4355 60954 4379 60956
rect 4435 60954 4459 60956
rect 4515 60954 4521 60956
rect 4275 60902 4277 60954
rect 4457 60902 4459 60954
rect 4213 60900 4219 60902
rect 4275 60900 4299 60902
rect 4355 60900 4379 60902
rect 4435 60900 4459 60902
rect 4515 60900 4521 60902
rect 4213 60880 4521 60900
rect 4213 59868 4521 59888
rect 4213 59866 4219 59868
rect 4275 59866 4299 59868
rect 4355 59866 4379 59868
rect 4435 59866 4459 59868
rect 4515 59866 4521 59868
rect 4275 59814 4277 59866
rect 4457 59814 4459 59866
rect 4213 59812 4219 59814
rect 4275 59812 4299 59814
rect 4355 59812 4379 59814
rect 4435 59812 4459 59814
rect 4515 59812 4521 59814
rect 4213 59792 4521 59812
rect 4213 58780 4521 58800
rect 4213 58778 4219 58780
rect 4275 58778 4299 58780
rect 4355 58778 4379 58780
rect 4435 58778 4459 58780
rect 4515 58778 4521 58780
rect 4275 58726 4277 58778
rect 4457 58726 4459 58778
rect 4213 58724 4219 58726
rect 4275 58724 4299 58726
rect 4355 58724 4379 58726
rect 4435 58724 4459 58726
rect 4515 58724 4521 58726
rect 4213 58704 4521 58724
rect 4213 57692 4521 57712
rect 4213 57690 4219 57692
rect 4275 57690 4299 57692
rect 4355 57690 4379 57692
rect 4435 57690 4459 57692
rect 4515 57690 4521 57692
rect 4275 57638 4277 57690
rect 4457 57638 4459 57690
rect 4213 57636 4219 57638
rect 4275 57636 4299 57638
rect 4355 57636 4379 57638
rect 4435 57636 4459 57638
rect 4515 57636 4521 57638
rect 4213 57616 4521 57636
rect 4213 56604 4521 56624
rect 4213 56602 4219 56604
rect 4275 56602 4299 56604
rect 4355 56602 4379 56604
rect 4435 56602 4459 56604
rect 4515 56602 4521 56604
rect 4275 56550 4277 56602
rect 4457 56550 4459 56602
rect 4213 56548 4219 56550
rect 4275 56548 4299 56550
rect 4355 56548 4379 56550
rect 4435 56548 4459 56550
rect 4515 56548 4521 56550
rect 4213 56528 4521 56548
rect 4213 55516 4521 55536
rect 4213 55514 4219 55516
rect 4275 55514 4299 55516
rect 4355 55514 4379 55516
rect 4435 55514 4459 55516
rect 4515 55514 4521 55516
rect 4275 55462 4277 55514
rect 4457 55462 4459 55514
rect 4213 55460 4219 55462
rect 4275 55460 4299 55462
rect 4355 55460 4379 55462
rect 4435 55460 4459 55462
rect 4515 55460 4521 55462
rect 4213 55440 4521 55460
rect 4213 54428 4521 54448
rect 4213 54426 4219 54428
rect 4275 54426 4299 54428
rect 4355 54426 4379 54428
rect 4435 54426 4459 54428
rect 4515 54426 4521 54428
rect 4275 54374 4277 54426
rect 4457 54374 4459 54426
rect 4213 54372 4219 54374
rect 4275 54372 4299 54374
rect 4355 54372 4379 54374
rect 4435 54372 4459 54374
rect 4515 54372 4521 54374
rect 4213 54352 4521 54372
rect 4213 53340 4521 53360
rect 4213 53338 4219 53340
rect 4275 53338 4299 53340
rect 4355 53338 4379 53340
rect 4435 53338 4459 53340
rect 4515 53338 4521 53340
rect 4275 53286 4277 53338
rect 4457 53286 4459 53338
rect 4213 53284 4219 53286
rect 4275 53284 4299 53286
rect 4355 53284 4379 53286
rect 4435 53284 4459 53286
rect 4515 53284 4521 53286
rect 4213 53264 4521 53284
rect 4213 52252 4521 52272
rect 4213 52250 4219 52252
rect 4275 52250 4299 52252
rect 4355 52250 4379 52252
rect 4435 52250 4459 52252
rect 4515 52250 4521 52252
rect 4275 52198 4277 52250
rect 4457 52198 4459 52250
rect 4213 52196 4219 52198
rect 4275 52196 4299 52198
rect 4355 52196 4379 52198
rect 4435 52196 4459 52198
rect 4515 52196 4521 52198
rect 4213 52176 4521 52196
rect 4213 51164 4521 51184
rect 4213 51162 4219 51164
rect 4275 51162 4299 51164
rect 4355 51162 4379 51164
rect 4435 51162 4459 51164
rect 4515 51162 4521 51164
rect 4275 51110 4277 51162
rect 4457 51110 4459 51162
rect 4213 51108 4219 51110
rect 4275 51108 4299 51110
rect 4355 51108 4379 51110
rect 4435 51108 4459 51110
rect 4515 51108 4521 51110
rect 4213 51088 4521 51108
rect 4213 50076 4521 50096
rect 4213 50074 4219 50076
rect 4275 50074 4299 50076
rect 4355 50074 4379 50076
rect 4435 50074 4459 50076
rect 4515 50074 4521 50076
rect 4275 50022 4277 50074
rect 4457 50022 4459 50074
rect 4213 50020 4219 50022
rect 4275 50020 4299 50022
rect 4355 50020 4379 50022
rect 4435 50020 4459 50022
rect 4515 50020 4521 50022
rect 4213 50000 4521 50020
rect 4160 49904 4212 49910
rect 4158 49872 4160 49881
rect 4212 49872 4214 49881
rect 4158 49807 4214 49816
rect 4213 48988 4521 49008
rect 4213 48986 4219 48988
rect 4275 48986 4299 48988
rect 4355 48986 4379 48988
rect 4435 48986 4459 48988
rect 4515 48986 4521 48988
rect 4275 48934 4277 48986
rect 4457 48934 4459 48986
rect 4213 48932 4219 48934
rect 4275 48932 4299 48934
rect 4355 48932 4379 48934
rect 4435 48932 4459 48934
rect 4515 48932 4521 48934
rect 4213 48912 4521 48932
rect 4632 48346 4660 74666
rect 5845 74556 6153 74576
rect 5845 74554 5851 74556
rect 5907 74554 5931 74556
rect 5987 74554 6011 74556
rect 6067 74554 6091 74556
rect 6147 74554 6153 74556
rect 5907 74502 5909 74554
rect 6089 74502 6091 74554
rect 5845 74500 5851 74502
rect 5907 74500 5931 74502
rect 5987 74500 6011 74502
rect 6067 74500 6091 74502
rect 6147 74500 6153 74502
rect 5845 74480 6153 74500
rect 4896 74384 4948 74390
rect 4896 74326 4948 74332
rect 4712 57928 4764 57934
rect 4712 57870 4764 57876
rect 4620 48340 4672 48346
rect 4620 48282 4672 48288
rect 4213 47900 4521 47920
rect 4213 47898 4219 47900
rect 4275 47898 4299 47900
rect 4355 47898 4379 47900
rect 4435 47898 4459 47900
rect 4515 47898 4521 47900
rect 4275 47846 4277 47898
rect 4457 47846 4459 47898
rect 4213 47844 4219 47846
rect 4275 47844 4299 47846
rect 4355 47844 4379 47846
rect 4435 47844 4459 47846
rect 4515 47844 4521 47846
rect 4213 47824 4521 47844
rect 4620 47184 4672 47190
rect 4620 47126 4672 47132
rect 4213 46812 4521 46832
rect 4213 46810 4219 46812
rect 4275 46810 4299 46812
rect 4355 46810 4379 46812
rect 4435 46810 4459 46812
rect 4515 46810 4521 46812
rect 4275 46758 4277 46810
rect 4457 46758 4459 46810
rect 4213 46756 4219 46758
rect 4275 46756 4299 46758
rect 4355 46756 4379 46758
rect 4435 46756 4459 46758
rect 4515 46756 4521 46758
rect 4213 46736 4521 46756
rect 4632 46458 4660 47126
rect 4540 46430 4660 46458
rect 4724 46442 4752 57870
rect 4908 51074 4936 74326
rect 5540 73636 5592 73642
rect 5540 73578 5592 73584
rect 5356 67108 5408 67114
rect 5356 67050 5408 67056
rect 5080 63980 5132 63986
rect 5080 63922 5132 63928
rect 4988 62892 5040 62898
rect 4988 62834 5040 62840
rect 4816 51046 4936 51074
rect 4816 49609 4844 51046
rect 4896 49904 4948 49910
rect 4896 49846 4948 49852
rect 4802 49600 4858 49609
rect 4802 49535 4858 49544
rect 4804 49428 4856 49434
rect 4804 49370 4856 49376
rect 4816 47190 4844 49370
rect 4804 47184 4856 47190
rect 4804 47126 4856 47132
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 4712 46436 4764 46442
rect 4540 45898 4568 46430
rect 4712 46378 4764 46384
rect 4620 46368 4672 46374
rect 4620 46310 4672 46316
rect 4528 45892 4580 45898
rect 4528 45834 4580 45840
rect 4213 45724 4521 45744
rect 4213 45722 4219 45724
rect 4275 45722 4299 45724
rect 4355 45722 4379 45724
rect 4435 45722 4459 45724
rect 4515 45722 4521 45724
rect 4275 45670 4277 45722
rect 4457 45670 4459 45722
rect 4213 45668 4219 45670
rect 4275 45668 4299 45670
rect 4355 45668 4379 45670
rect 4435 45668 4459 45670
rect 4515 45668 4521 45670
rect 4213 45648 4521 45668
rect 4213 44636 4521 44656
rect 4213 44634 4219 44636
rect 4275 44634 4299 44636
rect 4355 44634 4379 44636
rect 4435 44634 4459 44636
rect 4515 44634 4521 44636
rect 4275 44582 4277 44634
rect 4457 44582 4459 44634
rect 4213 44580 4219 44582
rect 4275 44580 4299 44582
rect 4355 44580 4379 44582
rect 4435 44580 4459 44582
rect 4515 44580 4521 44582
rect 4213 44560 4521 44580
rect 4436 44396 4488 44402
rect 4436 44338 4488 44344
rect 4448 44266 4476 44338
rect 4436 44260 4488 44266
rect 4436 44202 4488 44208
rect 4448 43926 4476 44202
rect 4436 43920 4488 43926
rect 4436 43862 4488 43868
rect 4213 43548 4521 43568
rect 4213 43546 4219 43548
rect 4275 43546 4299 43548
rect 4355 43546 4379 43548
rect 4435 43546 4459 43548
rect 4515 43546 4521 43548
rect 4275 43494 4277 43546
rect 4457 43494 4459 43546
rect 4213 43492 4219 43494
rect 4275 43492 4299 43494
rect 4355 43492 4379 43494
rect 4435 43492 4459 43494
rect 4515 43492 4521 43494
rect 4213 43472 4521 43492
rect 4526 43344 4582 43353
rect 4526 43279 4582 43288
rect 4540 42838 4568 43279
rect 4528 42832 4580 42838
rect 4528 42774 4580 42780
rect 4213 42460 4521 42480
rect 4213 42458 4219 42460
rect 4275 42458 4299 42460
rect 4355 42458 4379 42460
rect 4435 42458 4459 42460
rect 4515 42458 4521 42460
rect 4275 42406 4277 42458
rect 4457 42406 4459 42458
rect 4213 42404 4219 42406
rect 4275 42404 4299 42406
rect 4355 42404 4379 42406
rect 4435 42404 4459 42406
rect 4515 42404 4521 42406
rect 4213 42384 4521 42404
rect 4344 42288 4396 42294
rect 4158 42256 4214 42265
rect 4344 42230 4396 42236
rect 4158 42191 4214 42200
rect 4172 41682 4200 42191
rect 4160 41676 4212 41682
rect 4160 41618 4212 41624
rect 4356 41614 4384 42230
rect 4528 42220 4580 42226
rect 4528 42162 4580 42168
rect 4344 41608 4396 41614
rect 4344 41550 4396 41556
rect 4540 41528 4568 42162
rect 4632 41682 4660 46310
rect 4712 46096 4764 46102
rect 4712 46038 4764 46044
rect 4620 41676 4672 41682
rect 4620 41618 4672 41624
rect 4540 41500 4660 41528
rect 4213 41372 4521 41392
rect 4213 41370 4219 41372
rect 4275 41370 4299 41372
rect 4355 41370 4379 41372
rect 4435 41370 4459 41372
rect 4515 41370 4521 41372
rect 4275 41318 4277 41370
rect 4457 41318 4459 41370
rect 4213 41316 4219 41318
rect 4275 41316 4299 41318
rect 4355 41316 4379 41318
rect 4435 41316 4459 41318
rect 4515 41316 4521 41318
rect 4213 41296 4521 41316
rect 4213 40284 4521 40304
rect 4213 40282 4219 40284
rect 4275 40282 4299 40284
rect 4355 40282 4379 40284
rect 4435 40282 4459 40284
rect 4515 40282 4521 40284
rect 4275 40230 4277 40282
rect 4457 40230 4459 40282
rect 4213 40228 4219 40230
rect 4275 40228 4299 40230
rect 4355 40228 4379 40230
rect 4435 40228 4459 40230
rect 4515 40228 4521 40230
rect 4213 40208 4521 40228
rect 3976 40054 4028 40060
rect 4066 40080 4122 40089
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 3804 39302 3832 39986
rect 3884 39840 3936 39846
rect 3884 39782 3936 39788
rect 3896 39545 3924 39782
rect 3882 39536 3938 39545
rect 3882 39471 3938 39480
rect 3884 39432 3936 39438
rect 3884 39374 3936 39380
rect 3792 39296 3844 39302
rect 3792 39238 3844 39244
rect 3700 39024 3752 39030
rect 3700 38966 3752 38972
rect 3608 38820 3660 38826
rect 3608 38762 3660 38768
rect 3516 38480 3568 38486
rect 3516 38422 3568 38428
rect 3516 38344 3568 38350
rect 3516 38286 3568 38292
rect 3424 37256 3476 37262
rect 3424 37198 3476 37204
rect 3528 37074 3556 38286
rect 3436 37046 3556 37074
rect 3436 36310 3464 37046
rect 3514 36952 3570 36961
rect 3514 36887 3570 36896
rect 3528 36786 3556 36887
rect 3516 36780 3568 36786
rect 3516 36722 3568 36728
rect 3528 36689 3556 36722
rect 3514 36680 3570 36689
rect 3514 36615 3570 36624
rect 3424 36304 3476 36310
rect 3424 36246 3476 36252
rect 3516 36168 3568 36174
rect 3516 36110 3568 36116
rect 3528 35766 3556 36110
rect 3516 35760 3568 35766
rect 3516 35702 3568 35708
rect 3424 35080 3476 35086
rect 3424 35022 3476 35028
rect 3332 33992 3384 33998
rect 3332 33934 3384 33940
rect 3436 33930 3464 35022
rect 3424 33924 3476 33930
rect 3424 33866 3476 33872
rect 3330 33824 3386 33833
rect 3330 33759 3386 33768
rect 3240 29504 3292 29510
rect 3240 29446 3292 29452
rect 3252 25430 3280 29446
rect 3240 25424 3292 25430
rect 3240 25366 3292 25372
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3252 24721 3280 25230
rect 3344 24886 3372 33759
rect 3436 33522 3464 33866
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3436 32434 3464 33458
rect 3424 32428 3476 32434
rect 3424 32370 3476 32376
rect 3424 31816 3476 31822
rect 3424 31758 3476 31764
rect 3436 29306 3464 31758
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28529 3464 28902
rect 3422 28520 3478 28529
rect 3422 28455 3478 28464
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 3436 27305 3464 28018
rect 3422 27296 3478 27305
rect 3422 27231 3478 27240
rect 3528 27130 3556 35702
rect 3620 35698 3648 38762
rect 3608 35692 3660 35698
rect 3608 35634 3660 35640
rect 3712 35578 3740 38966
rect 3792 38956 3844 38962
rect 3792 38898 3844 38904
rect 3804 36786 3832 38898
rect 3896 36961 3924 39374
rect 3988 38962 4016 40054
rect 4066 40015 4122 40024
rect 4528 40044 4580 40050
rect 4528 39986 4580 39992
rect 4344 39840 4396 39846
rect 4344 39782 4396 39788
rect 4356 39506 4384 39782
rect 4344 39500 4396 39506
rect 4344 39442 4396 39448
rect 4068 39432 4120 39438
rect 4068 39374 4120 39380
rect 4080 39098 4108 39374
rect 4540 39370 4568 39986
rect 4528 39364 4580 39370
rect 4528 39306 4580 39312
rect 4213 39196 4521 39216
rect 4213 39194 4219 39196
rect 4275 39194 4299 39196
rect 4355 39194 4379 39196
rect 4435 39194 4459 39196
rect 4515 39194 4521 39196
rect 4275 39142 4277 39194
rect 4457 39142 4459 39194
rect 4213 39140 4219 39142
rect 4275 39140 4299 39142
rect 4355 39140 4379 39142
rect 4435 39140 4459 39142
rect 4515 39140 4521 39142
rect 4213 39120 4521 39140
rect 4068 39092 4120 39098
rect 4068 39034 4120 39040
rect 4066 38992 4122 39001
rect 3976 38956 4028 38962
rect 4066 38927 4068 38936
rect 3976 38898 4028 38904
rect 4120 38927 4122 38936
rect 4436 38956 4488 38962
rect 4068 38898 4120 38904
rect 4436 38898 4488 38904
rect 4080 38842 4108 38898
rect 3988 38814 4108 38842
rect 4342 38856 4398 38865
rect 3988 37369 4016 38814
rect 4342 38791 4398 38800
rect 4356 38418 4384 38791
rect 4344 38412 4396 38418
rect 4344 38354 4396 38360
rect 4448 38350 4476 38898
rect 4436 38344 4488 38350
rect 4436 38286 4488 38292
rect 4068 38208 4120 38214
rect 4068 38150 4120 38156
rect 3974 37360 4030 37369
rect 3974 37295 4030 37304
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3882 36952 3938 36961
rect 3882 36887 3938 36896
rect 3792 36780 3844 36786
rect 3844 36740 3924 36768
rect 3792 36722 3844 36728
rect 3792 36304 3844 36310
rect 3792 36246 3844 36252
rect 3620 35550 3740 35578
rect 3620 31754 3648 35550
rect 3698 35456 3754 35465
rect 3698 35391 3754 35400
rect 3608 31748 3660 31754
rect 3608 31690 3660 31696
rect 3606 31648 3662 31657
rect 3606 31583 3662 31592
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 3620 26874 3648 31583
rect 3712 29510 3740 35391
rect 3700 29504 3752 29510
rect 3700 29446 3752 29452
rect 3804 29288 3832 36246
rect 3896 36174 3924 36740
rect 3988 36378 4016 37198
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 3884 36168 3936 36174
rect 3884 36110 3936 36116
rect 4080 36020 4108 38150
rect 4213 38108 4521 38128
rect 4213 38106 4219 38108
rect 4275 38106 4299 38108
rect 4355 38106 4379 38108
rect 4435 38106 4459 38108
rect 4515 38106 4521 38108
rect 4275 38054 4277 38106
rect 4457 38054 4459 38106
rect 4213 38052 4219 38054
rect 4275 38052 4299 38054
rect 4355 38052 4379 38054
rect 4435 38052 4459 38054
rect 4515 38052 4521 38054
rect 4213 38032 4521 38052
rect 4213 37020 4521 37040
rect 4213 37018 4219 37020
rect 4275 37018 4299 37020
rect 4355 37018 4379 37020
rect 4435 37018 4459 37020
rect 4515 37018 4521 37020
rect 4275 36966 4277 37018
rect 4457 36966 4459 37018
rect 4213 36964 4219 36966
rect 4275 36964 4299 36966
rect 4355 36964 4379 36966
rect 4435 36964 4459 36966
rect 4515 36964 4521 36966
rect 4213 36944 4521 36964
rect 3712 29260 3832 29288
rect 3896 35992 4108 36020
rect 3712 27010 3740 29260
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 3804 28665 3832 29106
rect 3790 28656 3846 28665
rect 3790 28591 3846 28600
rect 3792 27668 3844 27674
rect 3792 27610 3844 27616
rect 3804 27470 3832 27610
rect 3792 27464 3844 27470
rect 3792 27406 3844 27412
rect 3712 26982 3832 27010
rect 3700 26920 3752 26926
rect 3436 26846 3648 26874
rect 3698 26888 3700 26897
rect 3752 26888 3754 26897
rect 3332 24880 3384 24886
rect 3332 24822 3384 24828
rect 3238 24712 3294 24721
rect 3238 24647 3294 24656
rect 3160 24262 3280 24290
rect 3148 24200 3200 24206
rect 3148 24142 3200 24148
rect 3160 23769 3188 24142
rect 3146 23760 3202 23769
rect 3146 23695 3202 23704
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 3160 22545 3188 22578
rect 3146 22536 3202 22545
rect 3146 22471 3202 22480
rect 3252 21468 3280 24262
rect 3344 21622 3372 24822
rect 3436 22098 3464 26846
rect 3698 26823 3754 26832
rect 3608 26784 3660 26790
rect 3606 26752 3608 26761
rect 3660 26752 3662 26761
rect 3606 26687 3662 26696
rect 3516 26376 3568 26382
rect 3514 26344 3516 26353
rect 3568 26344 3570 26353
rect 3514 26279 3570 26288
rect 3516 25424 3568 25430
rect 3516 25366 3568 25372
rect 3528 23254 3556 25366
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3516 23112 3568 23118
rect 3516 23054 3568 23060
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 3252 21440 3372 21468
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 3068 19514 3096 20538
rect 3160 19854 3188 21286
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3252 19922 3280 20198
rect 3240 19916 3292 19922
rect 3240 19858 3292 19864
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3056 19372 3108 19378
rect 3056 19314 3108 19320
rect 3068 19281 3096 19314
rect 3054 19272 3110 19281
rect 3054 19207 3110 19216
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3252 18601 3280 18702
rect 3238 18592 3294 18601
rect 3238 18527 3294 18536
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2608 17270 2636 17478
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 17105 2912 17138
rect 2870 17096 2926 17105
rect 2870 17031 2926 17040
rect 2582 16892 2890 16912
rect 2582 16890 2588 16892
rect 2644 16890 2668 16892
rect 2724 16890 2748 16892
rect 2804 16890 2828 16892
rect 2884 16890 2890 16892
rect 2644 16838 2646 16890
rect 2826 16838 2828 16890
rect 2582 16836 2588 16838
rect 2644 16836 2668 16838
rect 2724 16836 2748 16838
rect 2804 16836 2828 16838
rect 2884 16836 2890 16838
rect 2582 16816 2890 16836
rect 2976 16658 3004 17478
rect 3068 17377 3096 18226
rect 3054 17368 3110 17377
rect 3054 17303 3110 17312
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2582 15804 2890 15824
rect 2582 15802 2588 15804
rect 2644 15802 2668 15804
rect 2724 15802 2748 15804
rect 2804 15802 2828 15804
rect 2884 15802 2890 15804
rect 2644 15750 2646 15802
rect 2826 15750 2828 15802
rect 2582 15748 2588 15750
rect 2644 15748 2668 15750
rect 2724 15748 2748 15750
rect 2804 15748 2828 15750
rect 2884 15748 2890 15750
rect 2582 15728 2890 15748
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2056 15422 2176 15450
rect 2240 15422 2636 15450
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1858 13016 1914 13025
rect 1858 12951 1914 12960
rect 2056 12850 2084 15422
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 14414 2176 14962
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1398 9143 1454 9152
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8401 1440 8434
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1780 7954 1808 9522
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1400 7880 1452 7886
rect 1306 7848 1362 7857
rect 1400 7822 1452 7828
rect 1306 7783 1362 7792
rect 1320 7410 1348 7783
rect 1412 7449 1440 7822
rect 1398 7440 1454 7449
rect 1308 7404 1360 7410
rect 1398 7375 1454 7384
rect 1308 7346 1360 7352
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6633 1900 6666
rect 1858 6624 1914 6633
rect 1858 6559 1914 6568
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 2056 5710 2084 6258
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 1216 5296 1268 5302
rect 1216 5238 1268 5244
rect 1228 4146 1256 5238
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1306 3224 1362 3233
rect 1306 3159 1362 3168
rect 1320 2446 1348 3159
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1412 2689 1440 2926
rect 1398 2680 1454 2689
rect 1596 2650 1624 4558
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1688 3534 1716 4490
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1688 2650 1716 3470
rect 2056 2922 2084 5646
rect 2148 3058 2176 13874
rect 2240 11762 2268 15422
rect 2608 15366 2636 15422
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 3194 2268 4082
rect 2332 3738 2360 14350
rect 2424 11218 2452 15302
rect 2778 15192 2834 15201
rect 2778 15127 2780 15136
rect 2832 15127 2834 15136
rect 2780 15098 2832 15104
rect 2582 14716 2890 14736
rect 2582 14714 2588 14716
rect 2644 14714 2668 14716
rect 2724 14714 2748 14716
rect 2804 14714 2828 14716
rect 2884 14714 2890 14716
rect 2644 14662 2646 14714
rect 2826 14662 2828 14714
rect 2582 14660 2588 14662
rect 2644 14660 2668 14662
rect 2724 14660 2748 14662
rect 2804 14660 2828 14662
rect 2884 14660 2890 14662
rect 2582 14640 2890 14660
rect 2582 13628 2890 13648
rect 2582 13626 2588 13628
rect 2644 13626 2668 13628
rect 2724 13626 2748 13628
rect 2804 13626 2828 13628
rect 2884 13626 2890 13628
rect 2644 13574 2646 13626
rect 2826 13574 2828 13626
rect 2582 13572 2588 13574
rect 2644 13572 2668 13574
rect 2724 13572 2748 13574
rect 2804 13572 2828 13574
rect 2884 13572 2890 13574
rect 2582 13552 2890 13572
rect 2976 13530 3004 16458
rect 3068 15706 3096 16458
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3056 15020 3108 15026
rect 3056 14962 3108 14968
rect 3068 14414 3096 14962
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 3068 14074 3096 14350
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2792 12866 2820 13398
rect 2964 12912 3016 12918
rect 2792 12838 2912 12866
rect 2964 12854 3016 12860
rect 2884 12782 2912 12838
rect 2780 12776 2832 12782
rect 2778 12744 2780 12753
rect 2872 12776 2924 12782
rect 2832 12744 2834 12753
rect 2872 12718 2924 12724
rect 2778 12679 2834 12688
rect 2582 12540 2890 12560
rect 2582 12538 2588 12540
rect 2644 12538 2668 12540
rect 2724 12538 2748 12540
rect 2804 12538 2828 12540
rect 2884 12538 2890 12540
rect 2644 12486 2646 12538
rect 2826 12486 2828 12538
rect 2582 12484 2588 12486
rect 2644 12484 2668 12486
rect 2724 12484 2748 12486
rect 2804 12484 2828 12486
rect 2884 12484 2890 12486
rect 2582 12464 2890 12484
rect 2582 11452 2890 11472
rect 2582 11450 2588 11452
rect 2644 11450 2668 11452
rect 2724 11450 2748 11452
rect 2804 11450 2828 11452
rect 2884 11450 2890 11452
rect 2644 11398 2646 11450
rect 2826 11398 2828 11450
rect 2582 11396 2588 11398
rect 2644 11396 2668 11398
rect 2724 11396 2748 11398
rect 2804 11396 2828 11398
rect 2884 11396 2890 11398
rect 2582 11376 2890 11396
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2884 10674 2912 11086
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2582 10364 2890 10384
rect 2582 10362 2588 10364
rect 2644 10362 2668 10364
rect 2724 10362 2748 10364
rect 2804 10362 2828 10364
rect 2884 10362 2890 10364
rect 2644 10310 2646 10362
rect 2826 10310 2828 10362
rect 2582 10308 2588 10310
rect 2644 10308 2668 10310
rect 2724 10308 2748 10310
rect 2804 10308 2828 10310
rect 2884 10308 2890 10310
rect 2582 10288 2890 10308
rect 2976 10198 3004 12854
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2792 9518 2820 10066
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2582 9276 2890 9296
rect 2582 9274 2588 9276
rect 2644 9274 2668 9276
rect 2724 9274 2748 9276
rect 2804 9274 2828 9276
rect 2884 9274 2890 9276
rect 2644 9222 2646 9274
rect 2826 9222 2828 9274
rect 2582 9220 2588 9222
rect 2644 9220 2668 9222
rect 2724 9220 2748 9222
rect 2804 9220 2828 9222
rect 2884 9220 2890 9222
rect 2582 9200 2890 9220
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 2582 8188 2890 8208
rect 2582 8186 2588 8188
rect 2644 8186 2668 8188
rect 2724 8186 2748 8188
rect 2804 8186 2828 8188
rect 2884 8186 2890 8188
rect 2644 8134 2646 8186
rect 2826 8134 2828 8186
rect 2582 8132 2588 8134
rect 2644 8132 2668 8134
rect 2724 8132 2748 8134
rect 2804 8132 2828 8134
rect 2884 8132 2890 8134
rect 2582 8112 2890 8132
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 7313 2820 7346
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2582 7100 2890 7120
rect 2582 7098 2588 7100
rect 2644 7098 2668 7100
rect 2724 7098 2748 7100
rect 2804 7098 2828 7100
rect 2884 7098 2890 7100
rect 2644 7046 2646 7098
rect 2826 7046 2828 7098
rect 2582 7044 2588 7046
rect 2644 7044 2668 7046
rect 2724 7044 2748 7046
rect 2804 7044 2828 7046
rect 2884 7044 2890 7046
rect 2582 7024 2890 7044
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2884 6662 2912 6734
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2582 6012 2890 6032
rect 2582 6010 2588 6012
rect 2644 6010 2668 6012
rect 2724 6010 2748 6012
rect 2804 6010 2828 6012
rect 2884 6010 2890 6012
rect 2644 5958 2646 6010
rect 2826 5958 2828 6010
rect 2582 5956 2588 5958
rect 2644 5956 2668 5958
rect 2724 5956 2748 5958
rect 2804 5956 2828 5958
rect 2884 5956 2890 5958
rect 2582 5936 2890 5956
rect 2976 5914 3004 8842
rect 3068 6866 3096 13874
rect 3160 13802 3188 16730
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3252 16017 3280 16050
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3252 15026 3280 15098
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3238 14920 3294 14929
rect 3238 14855 3294 14864
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3252 13462 3280 14855
rect 3344 13938 3372 21440
rect 3528 20806 3556 23054
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3516 20528 3568 20534
rect 3516 20470 3568 20476
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3436 19553 3464 20402
rect 3528 20058 3556 20470
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3422 19544 3478 19553
rect 3422 19479 3478 19488
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3436 15162 3464 19382
rect 3620 17882 3648 26687
rect 3804 23322 3832 26982
rect 3792 23316 3844 23322
rect 3792 23258 3844 23264
rect 3896 22794 3924 35992
rect 4213 35932 4521 35952
rect 4213 35930 4219 35932
rect 4275 35930 4299 35932
rect 4355 35930 4379 35932
rect 4435 35930 4459 35932
rect 4515 35930 4521 35932
rect 4275 35878 4277 35930
rect 4457 35878 4459 35930
rect 4213 35876 4219 35878
rect 4275 35876 4299 35878
rect 4355 35876 4379 35878
rect 4435 35876 4459 35878
rect 4515 35876 4521 35878
rect 4213 35856 4521 35876
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 4172 35086 4200 35566
rect 4160 35080 4212 35086
rect 4160 35022 4212 35028
rect 4213 34844 4521 34864
rect 4213 34842 4219 34844
rect 4275 34842 4299 34844
rect 4355 34842 4379 34844
rect 4435 34842 4459 34844
rect 4515 34842 4521 34844
rect 4275 34790 4277 34842
rect 4457 34790 4459 34842
rect 4213 34788 4219 34790
rect 4275 34788 4299 34790
rect 4355 34788 4379 34790
rect 4435 34788 4459 34790
rect 4515 34788 4521 34790
rect 4213 34768 4521 34788
rect 4213 33756 4521 33776
rect 4213 33754 4219 33756
rect 4275 33754 4299 33756
rect 4355 33754 4379 33756
rect 4435 33754 4459 33756
rect 4515 33754 4521 33756
rect 4275 33702 4277 33754
rect 4457 33702 4459 33754
rect 4213 33700 4219 33702
rect 4275 33700 4299 33702
rect 4355 33700 4379 33702
rect 4435 33700 4459 33702
rect 4515 33700 4521 33702
rect 4213 33680 4521 33700
rect 4213 32668 4521 32688
rect 4213 32666 4219 32668
rect 4275 32666 4299 32668
rect 4355 32666 4379 32668
rect 4435 32666 4459 32668
rect 4515 32666 4521 32668
rect 4275 32614 4277 32666
rect 4457 32614 4459 32666
rect 4213 32612 4219 32614
rect 4275 32612 4299 32614
rect 4355 32612 4379 32614
rect 4435 32612 4459 32614
rect 4515 32612 4521 32614
rect 4213 32592 4521 32612
rect 3976 32428 4028 32434
rect 3976 32370 4028 32376
rect 3988 31822 4016 32370
rect 3976 31816 4028 31822
rect 3976 31758 4028 31764
rect 4068 31816 4120 31822
rect 4068 31758 4120 31764
rect 3976 31680 4028 31686
rect 3976 31622 4028 31628
rect 3988 28642 4016 31622
rect 4080 29034 4108 31758
rect 4213 31580 4521 31600
rect 4213 31578 4219 31580
rect 4275 31578 4299 31580
rect 4355 31578 4379 31580
rect 4435 31578 4459 31580
rect 4515 31578 4521 31580
rect 4275 31526 4277 31578
rect 4457 31526 4459 31578
rect 4213 31524 4219 31526
rect 4275 31524 4299 31526
rect 4355 31524 4379 31526
rect 4435 31524 4459 31526
rect 4515 31524 4521 31526
rect 4213 31504 4521 31524
rect 4213 30492 4521 30512
rect 4213 30490 4219 30492
rect 4275 30490 4299 30492
rect 4355 30490 4379 30492
rect 4435 30490 4459 30492
rect 4515 30490 4521 30492
rect 4275 30438 4277 30490
rect 4457 30438 4459 30490
rect 4213 30436 4219 30438
rect 4275 30436 4299 30438
rect 4355 30436 4379 30438
rect 4435 30436 4459 30438
rect 4515 30436 4521 30438
rect 4213 30416 4521 30436
rect 4213 29404 4521 29424
rect 4213 29402 4219 29404
rect 4275 29402 4299 29404
rect 4355 29402 4379 29404
rect 4435 29402 4459 29404
rect 4515 29402 4521 29404
rect 4275 29350 4277 29402
rect 4457 29350 4459 29402
rect 4213 29348 4219 29350
rect 4275 29348 4299 29350
rect 4355 29348 4379 29350
rect 4435 29348 4459 29350
rect 4515 29348 4521 29350
rect 4213 29328 4521 29348
rect 4068 29028 4120 29034
rect 4068 28970 4120 28976
rect 4632 28762 4660 41500
rect 4620 28756 4672 28762
rect 4620 28698 4672 28704
rect 4724 28642 4752 46038
rect 4816 41721 4844 46990
rect 4908 46209 4936 49846
rect 4894 46200 4950 46209
rect 4894 46135 4950 46144
rect 4896 46028 4948 46034
rect 4896 45970 4948 45976
rect 4802 41712 4858 41721
rect 4802 41647 4858 41656
rect 4804 41608 4856 41614
rect 4804 41550 4856 41556
rect 4816 33114 4844 41550
rect 4908 39642 4936 45970
rect 5000 45121 5028 62834
rect 5092 48210 5120 63922
rect 5172 63912 5224 63918
rect 5172 63854 5224 63860
rect 5184 49434 5212 63854
rect 5264 53032 5316 53038
rect 5264 52974 5316 52980
rect 5172 49428 5224 49434
rect 5172 49370 5224 49376
rect 5172 49292 5224 49298
rect 5172 49234 5224 49240
rect 5080 48204 5132 48210
rect 5080 48146 5132 48152
rect 5184 46560 5212 49234
rect 5092 46532 5212 46560
rect 4986 45112 5042 45121
rect 4986 45047 5042 45056
rect 5092 44962 5120 46532
rect 5172 46436 5224 46442
rect 5172 46378 5224 46384
rect 5000 44934 5120 44962
rect 5000 42226 5028 44934
rect 5080 44872 5132 44878
rect 5080 44814 5132 44820
rect 5092 43790 5120 44814
rect 5080 43784 5132 43790
rect 5080 43726 5132 43732
rect 5092 42294 5120 43726
rect 5080 42288 5132 42294
rect 5080 42230 5132 42236
rect 4988 42220 5040 42226
rect 4988 42162 5040 42168
rect 5092 42106 5120 42230
rect 5000 42078 5120 42106
rect 4896 39636 4948 39642
rect 4896 39578 4948 39584
rect 4894 39536 4950 39545
rect 4894 39471 4950 39480
rect 4908 38842 4936 39471
rect 5000 38962 5028 42078
rect 5078 41984 5134 41993
rect 5078 41919 5134 41928
rect 4988 38956 5040 38962
rect 4988 38898 5040 38904
rect 4908 38814 5028 38842
rect 5000 38282 5028 38814
rect 4988 38276 5040 38282
rect 4988 38218 5040 38224
rect 4896 36712 4948 36718
rect 4896 36654 4948 36660
rect 4804 33108 4856 33114
rect 4804 33050 4856 33056
rect 4804 32972 4856 32978
rect 4804 32914 4856 32920
rect 3988 28614 4108 28642
rect 3976 28552 4028 28558
rect 3976 28494 4028 28500
rect 3988 27985 4016 28494
rect 3974 27976 4030 27985
rect 3974 27911 4030 27920
rect 3974 27568 4030 27577
rect 3974 27503 4030 27512
rect 3988 27470 4016 27503
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 4080 27282 4108 28614
rect 4632 28614 4752 28642
rect 4213 28316 4521 28336
rect 4213 28314 4219 28316
rect 4275 28314 4299 28316
rect 4355 28314 4379 28316
rect 4435 28314 4459 28316
rect 4515 28314 4521 28316
rect 4275 28262 4277 28314
rect 4457 28262 4459 28314
rect 4213 28260 4219 28262
rect 4275 28260 4299 28262
rect 4355 28260 4379 28262
rect 4435 28260 4459 28262
rect 4515 28260 4521 28262
rect 4213 28240 4521 28260
rect 4632 27946 4660 28614
rect 4712 28484 4764 28490
rect 4712 28426 4764 28432
rect 4620 27940 4672 27946
rect 4620 27882 4672 27888
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 3712 22766 3924 22794
rect 3988 27254 4108 27282
rect 3712 22094 3740 22766
rect 3792 22704 3844 22710
rect 3792 22646 3844 22652
rect 3804 22234 3832 22646
rect 3988 22438 4016 27254
rect 4213 27228 4521 27248
rect 4213 27226 4219 27228
rect 4275 27226 4299 27228
rect 4355 27226 4379 27228
rect 4435 27226 4459 27228
rect 4515 27226 4521 27228
rect 4275 27174 4277 27226
rect 4457 27174 4459 27226
rect 4213 27172 4219 27174
rect 4275 27172 4299 27174
rect 4355 27172 4379 27174
rect 4435 27172 4459 27174
rect 4515 27172 4521 27174
rect 4213 27152 4521 27172
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 3976 22432 4028 22438
rect 3976 22374 4028 22380
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3712 22066 3832 22094
rect 3700 20936 3752 20942
rect 3700 20878 3752 20884
rect 3712 20602 3740 20878
rect 3700 20596 3752 20602
rect 3700 20538 3752 20544
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3528 15042 3556 17682
rect 3606 15192 3662 15201
rect 3606 15127 3608 15136
rect 3660 15127 3662 15136
rect 3608 15098 3660 15104
rect 3436 15014 3556 15042
rect 3608 15020 3660 15026
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 3436 13870 3464 15014
rect 3608 14962 3660 14968
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3332 13796 3384 13802
rect 3332 13738 3384 13744
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12850 3188 13262
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3160 10198 3188 12650
rect 3148 10192 3200 10198
rect 3148 10134 3200 10140
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3160 8498 3188 9998
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3068 5778 3096 6598
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2582 4924 2890 4944
rect 2582 4922 2588 4924
rect 2644 4922 2668 4924
rect 2724 4922 2748 4924
rect 2804 4922 2828 4924
rect 2884 4922 2890 4924
rect 2644 4870 2646 4922
rect 2826 4870 2828 4922
rect 2582 4868 2588 4870
rect 2644 4868 2668 4870
rect 2724 4868 2748 4870
rect 2804 4868 2828 4870
rect 2884 4868 2890 4870
rect 2582 4848 2890 4868
rect 2976 4729 3004 5646
rect 2962 4720 3018 4729
rect 2962 4655 3018 4664
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2332 3618 2360 3674
rect 2332 3590 2452 3618
rect 2424 3534 2452 3590
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 2516 2650 2544 4082
rect 3068 3942 3096 5714
rect 3160 4826 3188 8434
rect 3252 7886 3280 13194
rect 3344 11914 3372 13738
rect 3424 13728 3476 13734
rect 3424 13670 3476 13676
rect 3436 12306 3464 13670
rect 3528 13394 3556 14826
rect 3620 14396 3648 14962
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14550 3740 14894
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3620 14368 3740 14396
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 12714 3556 13330
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3344 11886 3464 11914
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3344 8974 3372 11698
rect 3436 9450 3464 11886
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3528 9722 3556 11154
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3252 7478 3280 7822
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 3252 5234 3280 7414
rect 3344 5914 3372 8910
rect 3436 7410 3464 9114
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3436 6914 3464 7346
rect 3528 7342 3556 9658
rect 3620 7546 3648 13874
rect 3712 12434 3740 14368
rect 3804 13938 3832 22066
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21729 4016 21966
rect 3974 21720 4030 21729
rect 3974 21655 4030 21664
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 3896 20777 3924 21490
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3882 20768 3938 20777
rect 3882 20703 3938 20712
rect 3884 20392 3936 20398
rect 3988 20369 4016 20878
rect 4080 20602 4108 27066
rect 4632 26994 4660 27406
rect 4724 27130 4752 28426
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4620 26988 4672 26994
rect 4672 26948 4752 26976
rect 4620 26930 4672 26936
rect 4724 26314 4752 26948
rect 4712 26308 4764 26314
rect 4712 26250 4764 26256
rect 4213 26140 4521 26160
rect 4213 26138 4219 26140
rect 4275 26138 4299 26140
rect 4355 26138 4379 26140
rect 4435 26138 4459 26140
rect 4515 26138 4521 26140
rect 4275 26086 4277 26138
rect 4457 26086 4459 26138
rect 4213 26084 4219 26086
rect 4275 26084 4299 26086
rect 4355 26084 4379 26086
rect 4435 26084 4459 26086
rect 4515 26084 4521 26086
rect 4213 26064 4521 26084
rect 4213 25052 4521 25072
rect 4213 25050 4219 25052
rect 4275 25050 4299 25052
rect 4355 25050 4379 25052
rect 4435 25050 4459 25052
rect 4515 25050 4521 25052
rect 4275 24998 4277 25050
rect 4457 24998 4459 25050
rect 4213 24996 4219 24998
rect 4275 24996 4299 24998
rect 4355 24996 4379 24998
rect 4435 24996 4459 24998
rect 4515 24996 4521 24998
rect 4213 24976 4521 24996
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4213 23964 4521 23984
rect 4213 23962 4219 23964
rect 4275 23962 4299 23964
rect 4355 23962 4379 23964
rect 4435 23962 4459 23964
rect 4515 23962 4521 23964
rect 4275 23910 4277 23962
rect 4457 23910 4459 23962
rect 4213 23908 4219 23910
rect 4275 23908 4299 23910
rect 4355 23908 4379 23910
rect 4435 23908 4459 23910
rect 4515 23908 4521 23910
rect 4213 23888 4521 23908
rect 4213 22876 4521 22896
rect 4213 22874 4219 22876
rect 4275 22874 4299 22876
rect 4355 22874 4379 22876
rect 4435 22874 4459 22876
rect 4515 22874 4521 22876
rect 4275 22822 4277 22874
rect 4457 22822 4459 22874
rect 4213 22820 4219 22822
rect 4275 22820 4299 22822
rect 4355 22820 4379 22822
rect 4435 22820 4459 22822
rect 4515 22820 4521 22822
rect 4213 22800 4521 22820
rect 4213 21788 4521 21808
rect 4213 21786 4219 21788
rect 4275 21786 4299 21788
rect 4355 21786 4379 21788
rect 4435 21786 4459 21788
rect 4515 21786 4521 21788
rect 4275 21734 4277 21786
rect 4457 21734 4459 21786
rect 4213 21732 4219 21734
rect 4275 21732 4299 21734
rect 4355 21732 4379 21734
rect 4435 21732 4459 21734
rect 4515 21732 4521 21734
rect 4213 21712 4521 21732
rect 4213 20700 4521 20720
rect 4213 20698 4219 20700
rect 4275 20698 4299 20700
rect 4355 20698 4379 20700
rect 4435 20698 4459 20700
rect 4515 20698 4521 20700
rect 4275 20646 4277 20698
rect 4457 20646 4459 20698
rect 4213 20644 4219 20646
rect 4275 20644 4299 20646
rect 4355 20644 4379 20646
rect 4435 20644 4459 20646
rect 4515 20644 4521 20646
rect 4213 20624 4521 20644
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 3884 20334 3936 20340
rect 3974 20360 4030 20369
rect 3896 17610 3924 20334
rect 3974 20295 4030 20304
rect 4080 19961 4108 20402
rect 4066 19952 4122 19961
rect 4066 19887 4122 19896
rect 4632 19786 4660 24754
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4213 19612 4521 19632
rect 4213 19610 4219 19612
rect 4275 19610 4299 19612
rect 4355 19610 4379 19612
rect 4435 19610 4459 19612
rect 4515 19610 4521 19612
rect 4275 19558 4277 19610
rect 4457 19558 4459 19610
rect 4213 19556 4219 19558
rect 4275 19556 4299 19558
rect 4355 19556 4379 19558
rect 4435 19556 4459 19558
rect 4515 19556 4521 19558
rect 4213 19536 4521 19556
rect 4213 18524 4521 18544
rect 4213 18522 4219 18524
rect 4275 18522 4299 18524
rect 4355 18522 4379 18524
rect 4435 18522 4459 18524
rect 4515 18522 4521 18524
rect 4275 18470 4277 18522
rect 4457 18470 4459 18522
rect 4213 18468 4219 18470
rect 4275 18468 4299 18470
rect 4355 18468 4379 18470
rect 4435 18468 4459 18470
rect 4515 18468 4521 18470
rect 4213 18448 4521 18468
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3896 14929 3924 17546
rect 4213 17436 4521 17456
rect 4213 17434 4219 17436
rect 4275 17434 4299 17436
rect 4355 17434 4379 17436
rect 4435 17434 4459 17436
rect 4515 17434 4521 17436
rect 4275 17382 4277 17434
rect 4457 17382 4459 17434
rect 4213 17380 4219 17382
rect 4275 17380 4299 17382
rect 4355 17380 4379 17382
rect 4435 17380 4459 17382
rect 4515 17380 4521 17382
rect 4213 17360 4521 17380
rect 4213 16348 4521 16368
rect 4213 16346 4219 16348
rect 4275 16346 4299 16348
rect 4355 16346 4379 16348
rect 4435 16346 4459 16348
rect 4515 16346 4521 16348
rect 4275 16294 4277 16346
rect 4457 16294 4459 16346
rect 4213 16292 4219 16294
rect 4275 16292 4299 16294
rect 4355 16292 4379 16294
rect 4435 16292 4459 16294
rect 4515 16292 4521 16294
rect 4213 16272 4521 16292
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3882 14920 3938 14929
rect 3882 14855 3938 14864
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 3896 13870 3924 14758
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 13977 4016 14350
rect 3974 13968 4030 13977
rect 3974 13903 4030 13912
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 4080 13734 4108 15506
rect 4213 15260 4521 15280
rect 4213 15258 4219 15260
rect 4275 15258 4299 15260
rect 4355 15258 4379 15260
rect 4435 15258 4459 15260
rect 4515 15258 4521 15260
rect 4275 15206 4277 15258
rect 4457 15206 4459 15258
rect 4213 15204 4219 15206
rect 4275 15204 4299 15206
rect 4355 15204 4379 15206
rect 4435 15204 4459 15206
rect 4515 15204 4521 15206
rect 4213 15184 4521 15204
rect 4160 14408 4212 14414
rect 4158 14376 4160 14385
rect 4212 14376 4214 14385
rect 4158 14311 4214 14320
rect 4213 14172 4521 14192
rect 4213 14170 4219 14172
rect 4275 14170 4299 14172
rect 4355 14170 4379 14172
rect 4435 14170 4459 14172
rect 4515 14170 4521 14172
rect 4275 14118 4277 14170
rect 4457 14118 4459 14170
rect 4213 14116 4219 14118
rect 4275 14116 4299 14118
rect 4355 14116 4379 14118
rect 4435 14116 4459 14118
rect 4515 14116 4521 14118
rect 4213 14096 4521 14116
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4066 13424 4122 13433
rect 4172 13410 4200 13874
rect 4122 13382 4200 13410
rect 4066 13359 4122 13368
rect 4632 13326 4660 19722
rect 4724 19718 4752 26250
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4724 14482 4752 19654
rect 4712 14476 4764 14482
rect 4712 14418 4764 14424
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4213 13084 4521 13104
rect 4213 13082 4219 13084
rect 4275 13082 4299 13084
rect 4355 13082 4379 13084
rect 4435 13082 4459 13084
rect 4515 13082 4521 13084
rect 4275 13030 4277 13082
rect 4457 13030 4459 13082
rect 4213 13028 4219 13030
rect 4275 13028 4299 13030
rect 4355 13028 4379 13030
rect 4435 13028 4459 13030
rect 4515 13028 4521 13030
rect 4213 13008 4521 13028
rect 3712 12406 3832 12434
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3712 8498 3740 10610
rect 3804 9178 3832 12406
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11150 3924 12174
rect 4213 11996 4521 12016
rect 4213 11994 4219 11996
rect 4275 11994 4299 11996
rect 4355 11994 4379 11996
rect 4435 11994 4459 11996
rect 4515 11994 4521 11996
rect 4275 11942 4277 11994
rect 4457 11942 4459 11994
rect 4213 11940 4219 11942
rect 4275 11940 4299 11942
rect 4355 11940 4379 11942
rect 4435 11940 4459 11942
rect 4515 11940 4521 11942
rect 4213 11920 4521 11940
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8809 3832 8910
rect 3790 8800 3846 8809
rect 3790 8735 3846 8744
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 7002 3648 7142
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3896 6914 3924 11086
rect 4213 10908 4521 10928
rect 4213 10906 4219 10908
rect 4275 10906 4299 10908
rect 4355 10906 4379 10908
rect 4435 10906 4459 10908
rect 4515 10906 4521 10908
rect 4275 10854 4277 10906
rect 4457 10854 4459 10906
rect 4213 10852 4219 10854
rect 4275 10852 4299 10854
rect 4355 10852 4379 10854
rect 4435 10852 4459 10854
rect 4515 10852 4521 10854
rect 4213 10832 4521 10852
rect 4213 9820 4521 9840
rect 4213 9818 4219 9820
rect 4275 9818 4299 9820
rect 4355 9818 4379 9820
rect 4435 9818 4459 9820
rect 4515 9818 4521 9820
rect 4275 9766 4277 9818
rect 4457 9766 4459 9818
rect 4213 9764 4219 9766
rect 4275 9764 4299 9766
rect 4355 9764 4379 9766
rect 4435 9764 4459 9766
rect 4515 9764 4521 9766
rect 4213 9744 4521 9764
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 8838 4016 9454
rect 4080 8974 4108 9522
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 4080 8634 4108 8910
rect 4213 8732 4521 8752
rect 4213 8730 4219 8732
rect 4275 8730 4299 8732
rect 4355 8730 4379 8732
rect 4435 8730 4459 8732
rect 4515 8730 4521 8732
rect 4275 8678 4277 8730
rect 4457 8678 4459 8730
rect 4213 8676 4219 8678
rect 4275 8676 4299 8678
rect 4355 8676 4379 8678
rect 4435 8676 4459 8678
rect 4515 8676 4521 8678
rect 4213 8656 4521 8676
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3436 6886 3556 6914
rect 3896 6886 4016 6914
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3436 5817 3464 6258
rect 3422 5808 3478 5817
rect 3422 5743 3478 5752
rect 3528 5370 3556 6886
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 6225 3832 6734
rect 3988 6662 4016 6886
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4080 6458 4108 8434
rect 4816 7818 4844 32914
rect 4908 28966 4936 36654
rect 5000 35601 5028 38218
rect 5092 36582 5120 41919
rect 5184 39914 5212 46378
rect 5276 46102 5304 52974
rect 5264 46096 5316 46102
rect 5264 46038 5316 46044
rect 5264 44328 5316 44334
rect 5264 44270 5316 44276
rect 5172 39908 5224 39914
rect 5172 39850 5224 39856
rect 5170 39808 5226 39817
rect 5170 39743 5226 39752
rect 5184 39574 5212 39743
rect 5172 39568 5224 39574
rect 5172 39510 5224 39516
rect 5172 39296 5224 39302
rect 5172 39238 5224 39244
rect 5080 36576 5132 36582
rect 5080 36518 5132 36524
rect 5078 36408 5134 36417
rect 5184 36378 5212 39238
rect 5276 36417 5304 44270
rect 5368 41585 5396 67050
rect 5448 63572 5500 63578
rect 5448 63514 5500 63520
rect 5460 62762 5488 63514
rect 5448 62756 5500 62762
rect 5448 62698 5500 62704
rect 5448 62484 5500 62490
rect 5448 62426 5500 62432
rect 5460 60636 5488 62426
rect 5552 60761 5580 73578
rect 5845 73468 6153 73488
rect 5845 73466 5851 73468
rect 5907 73466 5931 73468
rect 5987 73466 6011 73468
rect 6067 73466 6091 73468
rect 6147 73466 6153 73468
rect 5907 73414 5909 73466
rect 6089 73414 6091 73466
rect 5845 73412 5851 73414
rect 5907 73412 5931 73414
rect 5987 73412 6011 73414
rect 6067 73412 6091 73414
rect 6147 73412 6153 73414
rect 5845 73392 6153 73412
rect 5845 72380 6153 72400
rect 5845 72378 5851 72380
rect 5907 72378 5931 72380
rect 5987 72378 6011 72380
rect 6067 72378 6091 72380
rect 6147 72378 6153 72380
rect 5907 72326 5909 72378
rect 6089 72326 6091 72378
rect 5845 72324 5851 72326
rect 5907 72324 5931 72326
rect 5987 72324 6011 72326
rect 6067 72324 6091 72326
rect 6147 72324 6153 72326
rect 5845 72304 6153 72324
rect 5845 71292 6153 71312
rect 5845 71290 5851 71292
rect 5907 71290 5931 71292
rect 5987 71290 6011 71292
rect 6067 71290 6091 71292
rect 6147 71290 6153 71292
rect 5907 71238 5909 71290
rect 6089 71238 6091 71290
rect 5845 71236 5851 71238
rect 5907 71236 5931 71238
rect 5987 71236 6011 71238
rect 6067 71236 6091 71238
rect 6147 71236 6153 71238
rect 5845 71216 6153 71236
rect 6380 70394 6408 75890
rect 9109 75644 9417 75664
rect 9109 75642 9115 75644
rect 9171 75642 9195 75644
rect 9251 75642 9275 75644
rect 9331 75642 9355 75644
rect 9411 75642 9417 75644
rect 9171 75590 9173 75642
rect 9353 75590 9355 75642
rect 9109 75588 9115 75590
rect 9171 75588 9195 75590
rect 9251 75588 9275 75590
rect 9331 75588 9355 75590
rect 9411 75588 9417 75590
rect 9109 75568 9417 75588
rect 7477 75100 7785 75120
rect 7477 75098 7483 75100
rect 7539 75098 7563 75100
rect 7619 75098 7643 75100
rect 7699 75098 7723 75100
rect 7779 75098 7785 75100
rect 7539 75046 7541 75098
rect 7721 75046 7723 75098
rect 7477 75044 7483 75046
rect 7539 75044 7563 75046
rect 7619 75044 7643 75046
rect 7699 75044 7723 75046
rect 7779 75044 7785 75046
rect 7477 75024 7785 75044
rect 9876 74934 9904 76774
rect 10152 76537 10180 76978
rect 10138 76528 10194 76537
rect 10138 76463 10194 76472
rect 10232 75880 10284 75886
rect 10232 75822 10284 75828
rect 9956 75744 10008 75750
rect 10244 75721 10272 75822
rect 9956 75686 10008 75692
rect 10230 75712 10286 75721
rect 9864 74928 9916 74934
rect 9864 74870 9916 74876
rect 9968 74798 9996 75686
rect 10230 75647 10286 75656
rect 10140 75336 10192 75342
rect 10140 75278 10192 75284
rect 10152 74905 10180 75278
rect 10138 74896 10194 74905
rect 10138 74831 10194 74840
rect 9956 74792 10008 74798
rect 9956 74734 10008 74740
rect 8300 74656 8352 74662
rect 8300 74598 8352 74604
rect 7477 74012 7785 74032
rect 7477 74010 7483 74012
rect 7539 74010 7563 74012
rect 7619 74010 7643 74012
rect 7699 74010 7723 74012
rect 7779 74010 7785 74012
rect 7539 73958 7541 74010
rect 7721 73958 7723 74010
rect 7477 73956 7483 73958
rect 7539 73956 7563 73958
rect 7619 73956 7643 73958
rect 7699 73956 7723 73958
rect 7779 73956 7785 73958
rect 7477 73936 7785 73956
rect 7477 72924 7785 72944
rect 7477 72922 7483 72924
rect 7539 72922 7563 72924
rect 7619 72922 7643 72924
rect 7699 72922 7723 72924
rect 7779 72922 7785 72924
rect 7539 72870 7541 72922
rect 7721 72870 7723 72922
rect 7477 72868 7483 72870
rect 7539 72868 7563 72870
rect 7619 72868 7643 72870
rect 7699 72868 7723 72870
rect 7779 72868 7785 72870
rect 7477 72848 7785 72868
rect 7477 71836 7785 71856
rect 7477 71834 7483 71836
rect 7539 71834 7563 71836
rect 7619 71834 7643 71836
rect 7699 71834 7723 71836
rect 7779 71834 7785 71836
rect 7539 71782 7541 71834
rect 7721 71782 7723 71834
rect 7477 71780 7483 71782
rect 7539 71780 7563 71782
rect 7619 71780 7643 71782
rect 7699 71780 7723 71782
rect 7779 71780 7785 71782
rect 7477 71760 7785 71780
rect 7477 70748 7785 70768
rect 7477 70746 7483 70748
rect 7539 70746 7563 70748
rect 7619 70746 7643 70748
rect 7699 70746 7723 70748
rect 7779 70746 7785 70748
rect 7539 70694 7541 70746
rect 7721 70694 7723 70746
rect 7477 70692 7483 70694
rect 7539 70692 7563 70694
rect 7619 70692 7643 70694
rect 7699 70692 7723 70694
rect 7779 70692 7785 70694
rect 7477 70672 7785 70692
rect 7012 70440 7064 70446
rect 6380 70366 6592 70394
rect 7012 70382 7064 70388
rect 5845 70204 6153 70224
rect 5845 70202 5851 70204
rect 5907 70202 5931 70204
rect 5987 70202 6011 70204
rect 6067 70202 6091 70204
rect 6147 70202 6153 70204
rect 5907 70150 5909 70202
rect 6089 70150 6091 70202
rect 5845 70148 5851 70150
rect 5907 70148 5931 70150
rect 5987 70148 6011 70150
rect 6067 70148 6091 70150
rect 6147 70148 6153 70150
rect 5845 70128 6153 70148
rect 5724 69488 5776 69494
rect 5722 69456 5724 69465
rect 5776 69456 5778 69465
rect 5722 69391 5778 69400
rect 5845 69116 6153 69136
rect 5845 69114 5851 69116
rect 5907 69114 5931 69116
rect 5987 69114 6011 69116
rect 6067 69114 6091 69116
rect 6147 69114 6153 69116
rect 5907 69062 5909 69114
rect 6089 69062 6091 69114
rect 5845 69060 5851 69062
rect 5907 69060 5931 69062
rect 5987 69060 6011 69062
rect 6067 69060 6091 69062
rect 6147 69060 6153 69062
rect 5845 69040 6153 69060
rect 5845 68028 6153 68048
rect 5845 68026 5851 68028
rect 5907 68026 5931 68028
rect 5987 68026 6011 68028
rect 6067 68026 6091 68028
rect 6147 68026 6153 68028
rect 5907 67974 5909 68026
rect 6089 67974 6091 68026
rect 5845 67972 5851 67974
rect 5907 67972 5931 67974
rect 5987 67972 6011 67974
rect 6067 67972 6091 67974
rect 6147 67972 6153 67974
rect 5845 67952 6153 67972
rect 5845 66940 6153 66960
rect 5845 66938 5851 66940
rect 5907 66938 5931 66940
rect 5987 66938 6011 66940
rect 6067 66938 6091 66940
rect 6147 66938 6153 66940
rect 5907 66886 5909 66938
rect 6089 66886 6091 66938
rect 5845 66884 5851 66886
rect 5907 66884 5931 66886
rect 5987 66884 6011 66886
rect 6067 66884 6091 66886
rect 6147 66884 6153 66886
rect 5845 66864 6153 66884
rect 5845 65852 6153 65872
rect 5845 65850 5851 65852
rect 5907 65850 5931 65852
rect 5987 65850 6011 65852
rect 6067 65850 6091 65852
rect 6147 65850 6153 65852
rect 5907 65798 5909 65850
rect 6089 65798 6091 65850
rect 5845 65796 5851 65798
rect 5907 65796 5931 65798
rect 5987 65796 6011 65798
rect 6067 65796 6091 65798
rect 6147 65796 6153 65798
rect 5845 65776 6153 65796
rect 5632 65544 5684 65550
rect 5632 65486 5684 65492
rect 5538 60752 5594 60761
rect 5538 60687 5594 60696
rect 5460 60608 5580 60636
rect 5448 57248 5500 57254
rect 5448 57190 5500 57196
rect 5460 46034 5488 57190
rect 5552 48929 5580 60608
rect 5644 49065 5672 65486
rect 5845 64764 6153 64784
rect 5845 64762 5851 64764
rect 5907 64762 5931 64764
rect 5987 64762 6011 64764
rect 6067 64762 6091 64764
rect 6147 64762 6153 64764
rect 5907 64710 5909 64762
rect 6089 64710 6091 64762
rect 5845 64708 5851 64710
rect 5907 64708 5931 64710
rect 5987 64708 6011 64710
rect 6067 64708 6091 64710
rect 6147 64708 6153 64710
rect 5845 64688 6153 64708
rect 6276 63776 6328 63782
rect 6276 63718 6328 63724
rect 5845 63676 6153 63696
rect 5845 63674 5851 63676
rect 5907 63674 5931 63676
rect 5987 63674 6011 63676
rect 6067 63674 6091 63676
rect 6147 63674 6153 63676
rect 5907 63622 5909 63674
rect 6089 63622 6091 63674
rect 5845 63620 5851 63622
rect 5907 63620 5931 63622
rect 5987 63620 6011 63622
rect 6067 63620 6091 63622
rect 6147 63620 6153 63622
rect 5845 63600 6153 63620
rect 5724 63368 5776 63374
rect 5724 63310 5776 63316
rect 5736 54194 5764 63310
rect 5845 62588 6153 62608
rect 5845 62586 5851 62588
rect 5907 62586 5931 62588
rect 5987 62586 6011 62588
rect 6067 62586 6091 62588
rect 6147 62586 6153 62588
rect 5907 62534 5909 62586
rect 6089 62534 6091 62586
rect 5845 62532 5851 62534
rect 5907 62532 5931 62534
rect 5987 62532 6011 62534
rect 6067 62532 6091 62534
rect 6147 62532 6153 62534
rect 5845 62512 6153 62532
rect 5845 61500 6153 61520
rect 5845 61498 5851 61500
rect 5907 61498 5931 61500
rect 5987 61498 6011 61500
rect 6067 61498 6091 61500
rect 6147 61498 6153 61500
rect 5907 61446 5909 61498
rect 6089 61446 6091 61498
rect 5845 61444 5851 61446
rect 5907 61444 5931 61446
rect 5987 61444 6011 61446
rect 6067 61444 6091 61446
rect 6147 61444 6153 61446
rect 5845 61424 6153 61444
rect 6182 60616 6238 60625
rect 6182 60551 6238 60560
rect 5845 60412 6153 60432
rect 5845 60410 5851 60412
rect 5907 60410 5931 60412
rect 5987 60410 6011 60412
rect 6067 60410 6091 60412
rect 6147 60410 6153 60412
rect 5907 60358 5909 60410
rect 6089 60358 6091 60410
rect 5845 60356 5851 60358
rect 5907 60356 5931 60358
rect 5987 60356 6011 60358
rect 6067 60356 6091 60358
rect 6147 60356 6153 60358
rect 5845 60336 6153 60356
rect 5845 59324 6153 59344
rect 5845 59322 5851 59324
rect 5907 59322 5931 59324
rect 5987 59322 6011 59324
rect 6067 59322 6091 59324
rect 6147 59322 6153 59324
rect 5907 59270 5909 59322
rect 6089 59270 6091 59322
rect 5845 59268 5851 59270
rect 5907 59268 5931 59270
rect 5987 59268 6011 59270
rect 6067 59268 6091 59270
rect 6147 59268 6153 59270
rect 5845 59248 6153 59268
rect 5845 58236 6153 58256
rect 5845 58234 5851 58236
rect 5907 58234 5931 58236
rect 5987 58234 6011 58236
rect 6067 58234 6091 58236
rect 6147 58234 6153 58236
rect 5907 58182 5909 58234
rect 6089 58182 6091 58234
rect 5845 58180 5851 58182
rect 5907 58180 5931 58182
rect 5987 58180 6011 58182
rect 6067 58180 6091 58182
rect 6147 58180 6153 58182
rect 5845 58160 6153 58180
rect 5845 57148 6153 57168
rect 5845 57146 5851 57148
rect 5907 57146 5931 57148
rect 5987 57146 6011 57148
rect 6067 57146 6091 57148
rect 6147 57146 6153 57148
rect 5907 57094 5909 57146
rect 6089 57094 6091 57146
rect 5845 57092 5851 57094
rect 5907 57092 5931 57094
rect 5987 57092 6011 57094
rect 6067 57092 6091 57094
rect 6147 57092 6153 57094
rect 5845 57072 6153 57092
rect 5845 56060 6153 56080
rect 5845 56058 5851 56060
rect 5907 56058 5931 56060
rect 5987 56058 6011 56060
rect 6067 56058 6091 56060
rect 6147 56058 6153 56060
rect 5907 56006 5909 56058
rect 6089 56006 6091 56058
rect 5845 56004 5851 56006
rect 5907 56004 5931 56006
rect 5987 56004 6011 56006
rect 6067 56004 6091 56006
rect 6147 56004 6153 56006
rect 5845 55984 6153 56004
rect 5845 54972 6153 54992
rect 5845 54970 5851 54972
rect 5907 54970 5931 54972
rect 5987 54970 6011 54972
rect 6067 54970 6091 54972
rect 6147 54970 6153 54972
rect 5907 54918 5909 54970
rect 6089 54918 6091 54970
rect 5845 54916 5851 54918
rect 5907 54916 5931 54918
rect 5987 54916 6011 54918
rect 6067 54916 6091 54918
rect 6147 54916 6153 54918
rect 5845 54896 6153 54916
rect 5724 54188 5776 54194
rect 5724 54130 5776 54136
rect 5845 53884 6153 53904
rect 5845 53882 5851 53884
rect 5907 53882 5931 53884
rect 5987 53882 6011 53884
rect 6067 53882 6091 53884
rect 6147 53882 6153 53884
rect 5907 53830 5909 53882
rect 6089 53830 6091 53882
rect 5845 53828 5851 53830
rect 5907 53828 5931 53830
rect 5987 53828 6011 53830
rect 6067 53828 6091 53830
rect 6147 53828 6153 53830
rect 5845 53808 6153 53828
rect 5845 52796 6153 52816
rect 5845 52794 5851 52796
rect 5907 52794 5931 52796
rect 5987 52794 6011 52796
rect 6067 52794 6091 52796
rect 6147 52794 6153 52796
rect 5907 52742 5909 52794
rect 6089 52742 6091 52794
rect 5845 52740 5851 52742
rect 5907 52740 5931 52742
rect 5987 52740 6011 52742
rect 6067 52740 6091 52742
rect 6147 52740 6153 52742
rect 5845 52720 6153 52740
rect 5845 51708 6153 51728
rect 5845 51706 5851 51708
rect 5907 51706 5931 51708
rect 5987 51706 6011 51708
rect 6067 51706 6091 51708
rect 6147 51706 6153 51708
rect 5907 51654 5909 51706
rect 6089 51654 6091 51706
rect 5845 51652 5851 51654
rect 5907 51652 5931 51654
rect 5987 51652 6011 51654
rect 6067 51652 6091 51654
rect 6147 51652 6153 51654
rect 5845 51632 6153 51652
rect 5845 50620 6153 50640
rect 5845 50618 5851 50620
rect 5907 50618 5931 50620
rect 5987 50618 6011 50620
rect 6067 50618 6091 50620
rect 6147 50618 6153 50620
rect 5907 50566 5909 50618
rect 6089 50566 6091 50618
rect 5845 50564 5851 50566
rect 5907 50564 5931 50566
rect 5987 50564 6011 50566
rect 6067 50564 6091 50566
rect 6147 50564 6153 50566
rect 5845 50544 6153 50564
rect 5845 49532 6153 49552
rect 5845 49530 5851 49532
rect 5907 49530 5931 49532
rect 5987 49530 6011 49532
rect 6067 49530 6091 49532
rect 6147 49530 6153 49532
rect 5907 49478 5909 49530
rect 6089 49478 6091 49530
rect 5845 49476 5851 49478
rect 5907 49476 5931 49478
rect 5987 49476 6011 49478
rect 6067 49476 6091 49478
rect 6147 49476 6153 49478
rect 5845 49456 6153 49476
rect 5630 49056 5686 49065
rect 5630 48991 5686 49000
rect 5538 48920 5594 48929
rect 5538 48855 5594 48864
rect 6196 48634 6224 60551
rect 6288 57974 6316 63718
rect 6288 57946 6408 57974
rect 6276 54188 6328 54194
rect 6276 54130 6328 54136
rect 6104 48618 6224 48634
rect 6092 48612 6224 48618
rect 6144 48606 6224 48612
rect 6092 48554 6144 48560
rect 5724 48544 5776 48550
rect 5630 48512 5686 48521
rect 5724 48486 5776 48492
rect 6184 48544 6236 48550
rect 6184 48486 6236 48492
rect 5630 48447 5686 48456
rect 5538 48342 5594 48351
rect 5538 48277 5594 48286
rect 5448 46028 5500 46034
rect 5448 45970 5500 45976
rect 5448 45892 5500 45898
rect 5448 45834 5500 45840
rect 5460 44198 5488 45834
rect 5448 44192 5500 44198
rect 5448 44134 5500 44140
rect 5448 43716 5500 43722
rect 5448 43658 5500 43664
rect 5460 43110 5488 43658
rect 5448 43104 5500 43110
rect 5448 43046 5500 43052
rect 5354 41576 5410 41585
rect 5354 41511 5410 41520
rect 5356 41472 5408 41478
rect 5356 41414 5408 41420
rect 5262 36408 5318 36417
rect 5078 36343 5134 36352
rect 5172 36372 5224 36378
rect 4986 35592 5042 35601
rect 4986 35527 5042 35536
rect 4988 35488 5040 35494
rect 4988 35430 5040 35436
rect 4896 28960 4948 28966
rect 4896 28902 4948 28908
rect 4896 28756 4948 28762
rect 4896 28698 4948 28704
rect 4908 25974 4936 28698
rect 4896 25968 4948 25974
rect 4896 25910 4948 25916
rect 5000 25498 5028 35430
rect 5092 33810 5120 36343
rect 5262 36343 5318 36352
rect 5172 36314 5224 36320
rect 5368 35494 5396 41414
rect 5460 36718 5488 43046
rect 5552 41138 5580 48277
rect 5644 41698 5672 48447
rect 5736 46102 5764 48486
rect 5845 48444 6153 48464
rect 5845 48442 5851 48444
rect 5907 48442 5931 48444
rect 5987 48442 6011 48444
rect 6067 48442 6091 48444
rect 6147 48442 6153 48444
rect 5907 48390 5909 48442
rect 6089 48390 6091 48442
rect 5845 48388 5851 48390
rect 5907 48388 5931 48390
rect 5987 48388 6011 48390
rect 6067 48388 6091 48390
rect 6147 48388 6153 48390
rect 5845 48368 6153 48388
rect 6196 47841 6224 48486
rect 6182 47832 6238 47841
rect 6182 47767 6238 47776
rect 6184 47728 6236 47734
rect 6184 47670 6236 47676
rect 5845 47356 6153 47376
rect 5845 47354 5851 47356
rect 5907 47354 5931 47356
rect 5987 47354 6011 47356
rect 6067 47354 6091 47356
rect 6147 47354 6153 47356
rect 5907 47302 5909 47354
rect 6089 47302 6091 47354
rect 5845 47300 5851 47302
rect 5907 47300 5931 47302
rect 5987 47300 6011 47302
rect 6067 47300 6091 47302
rect 6147 47300 6153 47302
rect 5845 47280 6153 47300
rect 5845 46268 6153 46288
rect 5845 46266 5851 46268
rect 5907 46266 5931 46268
rect 5987 46266 6011 46268
rect 6067 46266 6091 46268
rect 6147 46266 6153 46268
rect 5907 46214 5909 46266
rect 6089 46214 6091 46266
rect 5845 46212 5851 46214
rect 5907 46212 5931 46214
rect 5987 46212 6011 46214
rect 6067 46212 6091 46214
rect 6147 46212 6153 46214
rect 5845 46192 6153 46212
rect 5724 46096 5776 46102
rect 5724 46038 5776 46044
rect 5722 45928 5778 45937
rect 5722 45863 5778 45872
rect 5736 42362 5764 45863
rect 5845 45180 6153 45200
rect 5845 45178 5851 45180
rect 5907 45178 5931 45180
rect 5987 45178 6011 45180
rect 6067 45178 6091 45180
rect 6147 45178 6153 45180
rect 5907 45126 5909 45178
rect 6089 45126 6091 45178
rect 5845 45124 5851 45126
rect 5907 45124 5931 45126
rect 5987 45124 6011 45126
rect 6067 45124 6091 45126
rect 6147 45124 6153 45126
rect 5845 45104 6153 45124
rect 5845 44092 6153 44112
rect 5845 44090 5851 44092
rect 5907 44090 5931 44092
rect 5987 44090 6011 44092
rect 6067 44090 6091 44092
rect 6147 44090 6153 44092
rect 5907 44038 5909 44090
rect 6089 44038 6091 44090
rect 5845 44036 5851 44038
rect 5907 44036 5931 44038
rect 5987 44036 6011 44038
rect 6067 44036 6091 44038
rect 6147 44036 6153 44038
rect 5845 44016 6153 44036
rect 5845 43004 6153 43024
rect 5845 43002 5851 43004
rect 5907 43002 5931 43004
rect 5987 43002 6011 43004
rect 6067 43002 6091 43004
rect 6147 43002 6153 43004
rect 5907 42950 5909 43002
rect 6089 42950 6091 43002
rect 5845 42948 5851 42950
rect 5907 42948 5931 42950
rect 5987 42948 6011 42950
rect 6067 42948 6091 42950
rect 6147 42948 6153 42950
rect 5845 42928 6153 42948
rect 5724 42356 5776 42362
rect 5724 42298 5776 42304
rect 5845 41916 6153 41936
rect 5845 41914 5851 41916
rect 5907 41914 5931 41916
rect 5987 41914 6011 41916
rect 6067 41914 6091 41916
rect 6147 41914 6153 41916
rect 5907 41862 5909 41914
rect 6089 41862 6091 41914
rect 5845 41860 5851 41862
rect 5907 41860 5931 41862
rect 5987 41860 6011 41862
rect 6067 41860 6091 41862
rect 6147 41860 6153 41862
rect 5845 41840 6153 41860
rect 6196 41698 6224 47670
rect 5644 41670 5764 41698
rect 5632 41608 5684 41614
rect 5632 41550 5684 41556
rect 5736 41562 5764 41670
rect 6104 41670 6224 41698
rect 5540 41132 5592 41138
rect 5540 41074 5592 41080
rect 5540 40996 5592 41002
rect 5540 40938 5592 40944
rect 5552 36854 5580 40938
rect 5644 37942 5672 41550
rect 5736 41534 5856 41562
rect 5724 41472 5776 41478
rect 5724 41414 5776 41420
rect 5828 41414 5856 41534
rect 6104 41478 6132 41670
rect 6182 41576 6238 41585
rect 6182 41511 6238 41520
rect 6092 41472 6144 41478
rect 6092 41414 6144 41420
rect 5632 37936 5684 37942
rect 5632 37878 5684 37884
rect 5540 36848 5592 36854
rect 5540 36790 5592 36796
rect 5448 36712 5500 36718
rect 5448 36654 5500 36660
rect 5448 36576 5500 36582
rect 5448 36518 5500 36524
rect 5356 35488 5408 35494
rect 5356 35430 5408 35436
rect 5262 35184 5318 35193
rect 5262 35119 5318 35128
rect 5092 33782 5212 33810
rect 5080 28960 5132 28966
rect 5080 28902 5132 28908
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 5092 24410 5120 28902
rect 5184 24682 5212 33782
rect 5172 24676 5224 24682
rect 5172 24618 5224 24624
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 5276 21078 5304 35119
rect 5356 33856 5408 33862
rect 5356 33798 5408 33804
rect 5368 22778 5396 33798
rect 5460 28694 5488 36518
rect 5540 36372 5592 36378
rect 5540 36314 5592 36320
rect 5552 33862 5580 36314
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5448 28688 5500 28694
rect 5448 28630 5500 28636
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5264 21072 5316 21078
rect 5264 21014 5316 21020
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5000 15366 5028 16050
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4213 7644 4521 7664
rect 4213 7642 4219 7644
rect 4275 7642 4299 7644
rect 4355 7642 4379 7644
rect 4435 7642 4459 7644
rect 4515 7642 4521 7644
rect 4275 7590 4277 7642
rect 4457 7590 4459 7642
rect 4213 7588 4219 7590
rect 4275 7588 4299 7590
rect 4355 7588 4379 7590
rect 4435 7588 4459 7590
rect 4515 7588 4521 7590
rect 4213 7568 4521 7588
rect 4213 6556 4521 6576
rect 4213 6554 4219 6556
rect 4275 6554 4299 6556
rect 4355 6554 4379 6556
rect 4435 6554 4459 6556
rect 4515 6554 4521 6556
rect 4275 6502 4277 6554
rect 4457 6502 4459 6554
rect 4213 6500 4219 6502
rect 4275 6500 4299 6502
rect 4355 6500 4379 6502
rect 4435 6500 4459 6502
rect 4515 6500 4521 6502
rect 4213 6480 4521 6500
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3884 6248 3936 6254
rect 3790 6216 3846 6225
rect 3884 6190 3936 6196
rect 3790 6151 3846 6160
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4282 3280 4422
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2582 3836 2890 3856
rect 2582 3834 2588 3836
rect 2644 3834 2668 3836
rect 2724 3834 2748 3836
rect 2804 3834 2828 3836
rect 2884 3834 2890 3836
rect 2644 3782 2646 3834
rect 2826 3782 2828 3834
rect 2582 3780 2588 3782
rect 2644 3780 2668 3782
rect 2724 3780 2748 3782
rect 2804 3780 2828 3782
rect 2884 3780 2890 3782
rect 2582 3760 2890 3780
rect 2870 3632 2926 3641
rect 2870 3567 2926 3576
rect 2884 3058 2912 3567
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3344 2922 3372 5102
rect 3528 4146 3556 5170
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3528 3534 3556 4082
rect 3620 4049 3648 4082
rect 3606 4040 3662 4049
rect 3606 3975 3662 3984
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3792 3460 3844 3466
rect 3792 3402 3844 3408
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 2582 2748 2890 2768
rect 2582 2746 2588 2748
rect 2644 2746 2668 2748
rect 2724 2746 2748 2748
rect 2804 2746 2828 2748
rect 2884 2746 2890 2748
rect 2644 2694 2646 2746
rect 2826 2694 2828 2746
rect 2582 2692 2588 2694
rect 2644 2692 2668 2694
rect 2724 2692 2748 2694
rect 2804 2692 2828 2694
rect 2884 2692 2890 2694
rect 2582 2672 2890 2692
rect 1398 2615 1454 2624
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 2504 2644 2556 2650
rect 2504 2586 2556 2592
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 2792 649 2820 2382
rect 2884 1465 2912 2382
rect 3528 2281 3556 2994
rect 3514 2272 3570 2281
rect 3514 2207 3570 2216
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3620 1057 3648 2994
rect 3804 2650 3832 3402
rect 3896 2650 3924 6190
rect 4816 6118 4844 7754
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5273 4016 5646
rect 4213 5468 4521 5488
rect 4213 5466 4219 5468
rect 4275 5466 4299 5468
rect 4355 5466 4379 5468
rect 4435 5466 4459 5468
rect 4515 5466 4521 5468
rect 4275 5414 4277 5466
rect 4457 5414 4459 5466
rect 4213 5412 4219 5414
rect 4275 5412 4299 5414
rect 4355 5412 4379 5414
rect 4435 5412 4459 5414
rect 4515 5412 4521 5414
rect 4213 5392 4521 5412
rect 3974 5264 4030 5273
rect 3974 5199 4030 5208
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3988 4457 4016 4558
rect 3974 4448 4030 4457
rect 3974 4383 4030 4392
rect 4213 4380 4521 4400
rect 4213 4378 4219 4380
rect 4275 4378 4299 4380
rect 4355 4378 4379 4380
rect 4435 4378 4459 4380
rect 4515 4378 4521 4380
rect 4275 4326 4277 4378
rect 4457 4326 4459 4378
rect 4213 4324 4219 4326
rect 4275 4324 4299 4326
rect 4355 4324 4379 4326
rect 4435 4324 4459 4326
rect 4515 4324 4521 4326
rect 4213 4304 4521 4324
rect 5552 4078 5580 32846
rect 5736 27334 5764 41414
rect 5828 41386 5948 41414
rect 5920 41002 5948 41386
rect 5908 40996 5960 41002
rect 5908 40938 5960 40944
rect 5845 40828 6153 40848
rect 5845 40826 5851 40828
rect 5907 40826 5931 40828
rect 5987 40826 6011 40828
rect 6067 40826 6091 40828
rect 6147 40826 6153 40828
rect 5907 40774 5909 40826
rect 6089 40774 6091 40826
rect 5845 40772 5851 40774
rect 5907 40772 5931 40774
rect 5987 40772 6011 40774
rect 6067 40772 6091 40774
rect 6147 40772 6153 40774
rect 5845 40752 6153 40772
rect 5845 39740 6153 39760
rect 5845 39738 5851 39740
rect 5907 39738 5931 39740
rect 5987 39738 6011 39740
rect 6067 39738 6091 39740
rect 6147 39738 6153 39740
rect 5907 39686 5909 39738
rect 6089 39686 6091 39738
rect 5845 39684 5851 39686
rect 5907 39684 5931 39686
rect 5987 39684 6011 39686
rect 6067 39684 6091 39686
rect 6147 39684 6153 39686
rect 5845 39664 6153 39684
rect 5845 38652 6153 38672
rect 5845 38650 5851 38652
rect 5907 38650 5931 38652
rect 5987 38650 6011 38652
rect 6067 38650 6091 38652
rect 6147 38650 6153 38652
rect 5907 38598 5909 38650
rect 6089 38598 6091 38650
rect 5845 38596 5851 38598
rect 5907 38596 5931 38598
rect 5987 38596 6011 38598
rect 6067 38596 6091 38598
rect 6147 38596 6153 38598
rect 5845 38576 6153 38596
rect 5845 37564 6153 37584
rect 5845 37562 5851 37564
rect 5907 37562 5931 37564
rect 5987 37562 6011 37564
rect 6067 37562 6091 37564
rect 6147 37562 6153 37564
rect 5907 37510 5909 37562
rect 6089 37510 6091 37562
rect 5845 37508 5851 37510
rect 5907 37508 5931 37510
rect 5987 37508 6011 37510
rect 6067 37508 6091 37510
rect 6147 37508 6153 37510
rect 5845 37488 6153 37508
rect 5845 36476 6153 36496
rect 5845 36474 5851 36476
rect 5907 36474 5931 36476
rect 5987 36474 6011 36476
rect 6067 36474 6091 36476
rect 6147 36474 6153 36476
rect 5907 36422 5909 36474
rect 6089 36422 6091 36474
rect 5845 36420 5851 36422
rect 5907 36420 5931 36422
rect 5987 36420 6011 36422
rect 6067 36420 6091 36422
rect 6147 36420 6153 36422
rect 5845 36400 6153 36420
rect 5845 35388 6153 35408
rect 5845 35386 5851 35388
rect 5907 35386 5931 35388
rect 5987 35386 6011 35388
rect 6067 35386 6091 35388
rect 6147 35386 6153 35388
rect 5907 35334 5909 35386
rect 6089 35334 6091 35386
rect 5845 35332 5851 35334
rect 5907 35332 5931 35334
rect 5987 35332 6011 35334
rect 6067 35332 6091 35334
rect 6147 35332 6153 35334
rect 5845 35312 6153 35332
rect 5845 34300 6153 34320
rect 5845 34298 5851 34300
rect 5907 34298 5931 34300
rect 5987 34298 6011 34300
rect 6067 34298 6091 34300
rect 6147 34298 6153 34300
rect 5907 34246 5909 34298
rect 6089 34246 6091 34298
rect 5845 34244 5851 34246
rect 5907 34244 5931 34246
rect 5987 34244 6011 34246
rect 6067 34244 6091 34246
rect 6147 34244 6153 34246
rect 5845 34224 6153 34244
rect 5845 33212 6153 33232
rect 5845 33210 5851 33212
rect 5907 33210 5931 33212
rect 5987 33210 6011 33212
rect 6067 33210 6091 33212
rect 6147 33210 6153 33212
rect 5907 33158 5909 33210
rect 6089 33158 6091 33210
rect 5845 33156 5851 33158
rect 5907 33156 5931 33158
rect 5987 33156 6011 33158
rect 6067 33156 6091 33158
rect 6147 33156 6153 33158
rect 5845 33136 6153 33156
rect 5845 32124 6153 32144
rect 5845 32122 5851 32124
rect 5907 32122 5931 32124
rect 5987 32122 6011 32124
rect 6067 32122 6091 32124
rect 6147 32122 6153 32124
rect 5907 32070 5909 32122
rect 6089 32070 6091 32122
rect 5845 32068 5851 32070
rect 5907 32068 5931 32070
rect 5987 32068 6011 32070
rect 6067 32068 6091 32070
rect 6147 32068 6153 32070
rect 5845 32048 6153 32068
rect 5845 31036 6153 31056
rect 5845 31034 5851 31036
rect 5907 31034 5931 31036
rect 5987 31034 6011 31036
rect 6067 31034 6091 31036
rect 6147 31034 6153 31036
rect 5907 30982 5909 31034
rect 6089 30982 6091 31034
rect 5845 30980 5851 30982
rect 5907 30980 5931 30982
rect 5987 30980 6011 30982
rect 6067 30980 6091 30982
rect 6147 30980 6153 30982
rect 5845 30960 6153 30980
rect 5845 29948 6153 29968
rect 5845 29946 5851 29948
rect 5907 29946 5931 29948
rect 5987 29946 6011 29948
rect 6067 29946 6091 29948
rect 6147 29946 6153 29948
rect 5907 29894 5909 29946
rect 6089 29894 6091 29946
rect 5845 29892 5851 29894
rect 5907 29892 5931 29894
rect 5987 29892 6011 29894
rect 6067 29892 6091 29894
rect 6147 29892 6153 29894
rect 5845 29872 6153 29892
rect 5845 28860 6153 28880
rect 5845 28858 5851 28860
rect 5907 28858 5931 28860
rect 5987 28858 6011 28860
rect 6067 28858 6091 28860
rect 6147 28858 6153 28860
rect 5907 28806 5909 28858
rect 6089 28806 6091 28858
rect 5845 28804 5851 28806
rect 5907 28804 5931 28806
rect 5987 28804 6011 28806
rect 6067 28804 6091 28806
rect 6147 28804 6153 28806
rect 5845 28784 6153 28804
rect 5845 27772 6153 27792
rect 5845 27770 5851 27772
rect 5907 27770 5931 27772
rect 5987 27770 6011 27772
rect 6067 27770 6091 27772
rect 6147 27770 6153 27772
rect 5907 27718 5909 27770
rect 6089 27718 6091 27770
rect 5845 27716 5851 27718
rect 5907 27716 5931 27718
rect 5987 27716 6011 27718
rect 6067 27716 6091 27718
rect 6147 27716 6153 27718
rect 5845 27696 6153 27716
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5845 26684 6153 26704
rect 5845 26682 5851 26684
rect 5907 26682 5931 26684
rect 5987 26682 6011 26684
rect 6067 26682 6091 26684
rect 6147 26682 6153 26684
rect 5907 26630 5909 26682
rect 6089 26630 6091 26682
rect 5845 26628 5851 26630
rect 5907 26628 5931 26630
rect 5987 26628 6011 26630
rect 6067 26628 6091 26630
rect 6147 26628 6153 26630
rect 5845 26608 6153 26628
rect 5845 25596 6153 25616
rect 5845 25594 5851 25596
rect 5907 25594 5931 25596
rect 5987 25594 6011 25596
rect 6067 25594 6091 25596
rect 6147 25594 6153 25596
rect 5907 25542 5909 25594
rect 6089 25542 6091 25594
rect 5845 25540 5851 25542
rect 5907 25540 5931 25542
rect 5987 25540 6011 25542
rect 6067 25540 6091 25542
rect 6147 25540 6153 25542
rect 5845 25520 6153 25540
rect 5845 24508 6153 24528
rect 5845 24506 5851 24508
rect 5907 24506 5931 24508
rect 5987 24506 6011 24508
rect 6067 24506 6091 24508
rect 6147 24506 6153 24508
rect 5907 24454 5909 24506
rect 6089 24454 6091 24506
rect 5845 24452 5851 24454
rect 5907 24452 5931 24454
rect 5987 24452 6011 24454
rect 6067 24452 6091 24454
rect 6147 24452 6153 24454
rect 5845 24432 6153 24452
rect 5845 23420 6153 23440
rect 5845 23418 5851 23420
rect 5907 23418 5931 23420
rect 5987 23418 6011 23420
rect 6067 23418 6091 23420
rect 6147 23418 6153 23420
rect 5907 23366 5909 23418
rect 6089 23366 6091 23418
rect 5845 23364 5851 23366
rect 5907 23364 5931 23366
rect 5987 23364 6011 23366
rect 6067 23364 6091 23366
rect 6147 23364 6153 23366
rect 5845 23344 6153 23364
rect 5845 22332 6153 22352
rect 5845 22330 5851 22332
rect 5907 22330 5931 22332
rect 5987 22330 6011 22332
rect 6067 22330 6091 22332
rect 6147 22330 6153 22332
rect 5907 22278 5909 22330
rect 6089 22278 6091 22330
rect 5845 22276 5851 22278
rect 5907 22276 5931 22278
rect 5987 22276 6011 22278
rect 6067 22276 6091 22278
rect 6147 22276 6153 22278
rect 5845 22256 6153 22276
rect 5845 21244 6153 21264
rect 5845 21242 5851 21244
rect 5907 21242 5931 21244
rect 5987 21242 6011 21244
rect 6067 21242 6091 21244
rect 6147 21242 6153 21244
rect 5907 21190 5909 21242
rect 6089 21190 6091 21242
rect 5845 21188 5851 21190
rect 5907 21188 5931 21190
rect 5987 21188 6011 21190
rect 6067 21188 6091 21190
rect 6147 21188 6153 21190
rect 5845 21168 6153 21188
rect 5845 20156 6153 20176
rect 5845 20154 5851 20156
rect 5907 20154 5931 20156
rect 5987 20154 6011 20156
rect 6067 20154 6091 20156
rect 6147 20154 6153 20156
rect 5907 20102 5909 20154
rect 6089 20102 6091 20154
rect 5845 20100 5851 20102
rect 5907 20100 5931 20102
rect 5987 20100 6011 20102
rect 6067 20100 6091 20102
rect 6147 20100 6153 20102
rect 5845 20080 6153 20100
rect 5845 19068 6153 19088
rect 5845 19066 5851 19068
rect 5907 19066 5931 19068
rect 5987 19066 6011 19068
rect 6067 19066 6091 19068
rect 6147 19066 6153 19068
rect 5907 19014 5909 19066
rect 6089 19014 6091 19066
rect 5845 19012 5851 19014
rect 5907 19012 5931 19014
rect 5987 19012 6011 19014
rect 6067 19012 6091 19014
rect 6147 19012 6153 19014
rect 5845 18992 6153 19012
rect 5845 17980 6153 18000
rect 5845 17978 5851 17980
rect 5907 17978 5931 17980
rect 5987 17978 6011 17980
rect 6067 17978 6091 17980
rect 6147 17978 6153 17980
rect 5907 17926 5909 17978
rect 6089 17926 6091 17978
rect 5845 17924 5851 17926
rect 5907 17924 5931 17926
rect 5987 17924 6011 17926
rect 6067 17924 6091 17926
rect 6147 17924 6153 17926
rect 5845 17904 6153 17924
rect 5845 16892 6153 16912
rect 5845 16890 5851 16892
rect 5907 16890 5931 16892
rect 5987 16890 6011 16892
rect 6067 16890 6091 16892
rect 6147 16890 6153 16892
rect 5907 16838 5909 16890
rect 6089 16838 6091 16890
rect 5845 16836 5851 16838
rect 5907 16836 5931 16838
rect 5987 16836 6011 16838
rect 6067 16836 6091 16838
rect 6147 16836 6153 16838
rect 5845 16816 6153 16836
rect 5845 15804 6153 15824
rect 5845 15802 5851 15804
rect 5907 15802 5931 15804
rect 5987 15802 6011 15804
rect 6067 15802 6091 15804
rect 6147 15802 6153 15804
rect 5907 15750 5909 15802
rect 6089 15750 6091 15802
rect 5845 15748 5851 15750
rect 5907 15748 5931 15750
rect 5987 15748 6011 15750
rect 6067 15748 6091 15750
rect 6147 15748 6153 15750
rect 5845 15728 6153 15748
rect 5845 14716 6153 14736
rect 5845 14714 5851 14716
rect 5907 14714 5931 14716
rect 5987 14714 6011 14716
rect 6067 14714 6091 14716
rect 6147 14714 6153 14716
rect 5907 14662 5909 14714
rect 6089 14662 6091 14714
rect 5845 14660 5851 14662
rect 5907 14660 5931 14662
rect 5987 14660 6011 14662
rect 6067 14660 6091 14662
rect 6147 14660 6153 14662
rect 5845 14640 6153 14660
rect 5845 13628 6153 13648
rect 5845 13626 5851 13628
rect 5907 13626 5931 13628
rect 5987 13626 6011 13628
rect 6067 13626 6091 13628
rect 6147 13626 6153 13628
rect 5907 13574 5909 13626
rect 6089 13574 6091 13626
rect 5845 13572 5851 13574
rect 5907 13572 5931 13574
rect 5987 13572 6011 13574
rect 6067 13572 6091 13574
rect 6147 13572 6153 13574
rect 5845 13552 6153 13572
rect 5845 12540 6153 12560
rect 5845 12538 5851 12540
rect 5907 12538 5931 12540
rect 5987 12538 6011 12540
rect 6067 12538 6091 12540
rect 6147 12538 6153 12540
rect 5907 12486 5909 12538
rect 6089 12486 6091 12538
rect 5845 12484 5851 12486
rect 5907 12484 5931 12486
rect 5987 12484 6011 12486
rect 6067 12484 6091 12486
rect 6147 12484 6153 12486
rect 5845 12464 6153 12484
rect 6196 11898 6224 41511
rect 6288 41274 6316 54130
rect 6380 41614 6408 57946
rect 6564 49201 6592 70366
rect 6920 66564 6972 66570
rect 6920 66506 6972 66512
rect 6828 54664 6880 54670
rect 6828 54606 6880 54612
rect 6644 53168 6696 53174
rect 6644 53110 6696 53116
rect 6550 49192 6606 49201
rect 6550 49127 6606 49136
rect 6460 48884 6512 48890
rect 6460 48826 6512 48832
rect 6472 46481 6500 48826
rect 6458 46472 6514 46481
rect 6458 46407 6514 46416
rect 6656 46322 6684 53110
rect 6840 51074 6868 54606
rect 6472 46294 6684 46322
rect 6748 51046 6868 51074
rect 6368 41608 6420 41614
rect 6368 41550 6420 41556
rect 6472 41546 6500 46294
rect 6748 46186 6776 51046
rect 6826 48648 6882 48657
rect 6826 48583 6882 48592
rect 6564 46158 6776 46186
rect 6460 41540 6512 41546
rect 6460 41482 6512 41488
rect 6368 41472 6420 41478
rect 6368 41414 6420 41420
rect 6458 41440 6514 41449
rect 6276 41268 6328 41274
rect 6276 41210 6328 41216
rect 6276 41132 6328 41138
rect 6276 41074 6328 41080
rect 6288 35154 6316 41074
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 6274 27432 6330 27441
rect 6274 27367 6276 27376
rect 6328 27367 6330 27376
rect 6276 27338 6328 27344
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 5845 11452 6153 11472
rect 5845 11450 5851 11452
rect 5907 11450 5931 11452
rect 5987 11450 6011 11452
rect 6067 11450 6091 11452
rect 6147 11450 6153 11452
rect 5907 11398 5909 11450
rect 6089 11398 6091 11450
rect 5845 11396 5851 11398
rect 5907 11396 5931 11398
rect 5987 11396 6011 11398
rect 6067 11396 6091 11398
rect 6147 11396 6153 11398
rect 5845 11376 6153 11396
rect 5845 10364 6153 10384
rect 5845 10362 5851 10364
rect 5907 10362 5931 10364
rect 5987 10362 6011 10364
rect 6067 10362 6091 10364
rect 6147 10362 6153 10364
rect 5907 10310 5909 10362
rect 6089 10310 6091 10362
rect 5845 10308 5851 10310
rect 5907 10308 5931 10310
rect 5987 10308 6011 10310
rect 6067 10308 6091 10310
rect 6147 10308 6153 10310
rect 5845 10288 6153 10308
rect 5845 9276 6153 9296
rect 5845 9274 5851 9276
rect 5907 9274 5931 9276
rect 5987 9274 6011 9276
rect 6067 9274 6091 9276
rect 6147 9274 6153 9276
rect 5907 9222 5909 9274
rect 6089 9222 6091 9274
rect 5845 9220 5851 9222
rect 5907 9220 5931 9222
rect 5987 9220 6011 9222
rect 6067 9220 6091 9222
rect 6147 9220 6153 9222
rect 5845 9200 6153 9220
rect 5845 8188 6153 8208
rect 5845 8186 5851 8188
rect 5907 8186 5931 8188
rect 5987 8186 6011 8188
rect 6067 8186 6091 8188
rect 6147 8186 6153 8188
rect 5907 8134 5909 8186
rect 6089 8134 6091 8186
rect 5845 8132 5851 8134
rect 5907 8132 5931 8134
rect 5987 8132 6011 8134
rect 6067 8132 6091 8134
rect 6147 8132 6153 8134
rect 5845 8112 6153 8132
rect 5845 7100 6153 7120
rect 5845 7098 5851 7100
rect 5907 7098 5931 7100
rect 5987 7098 6011 7100
rect 6067 7098 6091 7100
rect 6147 7098 6153 7100
rect 5907 7046 5909 7098
rect 6089 7046 6091 7098
rect 5845 7044 5851 7046
rect 5907 7044 5931 7046
rect 5987 7044 6011 7046
rect 6067 7044 6091 7046
rect 6147 7044 6153 7046
rect 5845 7024 6153 7044
rect 6380 6914 6408 41414
rect 6458 41375 6514 41384
rect 6288 6886 6408 6914
rect 5845 6012 6153 6032
rect 5845 6010 5851 6012
rect 5907 6010 5931 6012
rect 5987 6010 6011 6012
rect 6067 6010 6091 6012
rect 6147 6010 6153 6012
rect 5907 5958 5909 6010
rect 6089 5958 6091 6010
rect 5845 5956 5851 5958
rect 5907 5956 5931 5958
rect 5987 5956 6011 5958
rect 6067 5956 6091 5958
rect 6147 5956 6153 5958
rect 5845 5936 6153 5956
rect 5845 4924 6153 4944
rect 5845 4922 5851 4924
rect 5907 4922 5931 4924
rect 5987 4922 6011 4924
rect 6067 4922 6091 4924
rect 6147 4922 6153 4924
rect 5907 4870 5909 4922
rect 6089 4870 6091 4922
rect 5845 4868 5851 4870
rect 5907 4868 5931 4870
rect 5987 4868 6011 4870
rect 6067 4868 6091 4870
rect 6147 4868 6153 4870
rect 5845 4848 6153 4868
rect 6288 4758 6316 6886
rect 6472 6730 6500 41375
rect 6564 32502 6592 46158
rect 6644 46096 6696 46102
rect 6644 46038 6696 46044
rect 6734 46064 6790 46073
rect 6552 32496 6604 32502
rect 6552 32438 6604 32444
rect 6656 10266 6684 46038
rect 6734 45999 6790 46008
rect 6748 41585 6776 45999
rect 6734 41576 6790 41585
rect 6734 41511 6790 41520
rect 6734 41304 6790 41313
rect 6734 41239 6790 41248
rect 6748 11286 6776 41239
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6840 5846 6868 48583
rect 6932 35834 6960 66506
rect 7024 46481 7052 70382
rect 7477 69660 7785 69680
rect 7477 69658 7483 69660
rect 7539 69658 7563 69660
rect 7619 69658 7643 69660
rect 7699 69658 7723 69660
rect 7779 69658 7785 69660
rect 7539 69606 7541 69658
rect 7721 69606 7723 69658
rect 7477 69604 7483 69606
rect 7539 69604 7563 69606
rect 7619 69604 7643 69606
rect 7699 69604 7723 69606
rect 7779 69604 7785 69606
rect 7477 69584 7785 69604
rect 7477 68572 7785 68592
rect 7477 68570 7483 68572
rect 7539 68570 7563 68572
rect 7619 68570 7643 68572
rect 7699 68570 7723 68572
rect 7779 68570 7785 68572
rect 7539 68518 7541 68570
rect 7721 68518 7723 68570
rect 7477 68516 7483 68518
rect 7539 68516 7563 68518
rect 7619 68516 7643 68518
rect 7699 68516 7723 68518
rect 7779 68516 7785 68518
rect 7477 68496 7785 68516
rect 7104 68264 7156 68270
rect 7104 68206 7156 68212
rect 7010 46472 7066 46481
rect 7010 46407 7066 46416
rect 7116 46322 7144 68206
rect 7477 67484 7785 67504
rect 7477 67482 7483 67484
rect 7539 67482 7563 67484
rect 7619 67482 7643 67484
rect 7699 67482 7723 67484
rect 7779 67482 7785 67484
rect 7539 67430 7541 67482
rect 7721 67430 7723 67482
rect 7477 67428 7483 67430
rect 7539 67428 7563 67430
rect 7619 67428 7643 67430
rect 7699 67428 7723 67430
rect 7779 67428 7785 67430
rect 7477 67408 7785 67428
rect 7477 66396 7785 66416
rect 7477 66394 7483 66396
rect 7539 66394 7563 66396
rect 7619 66394 7643 66396
rect 7699 66394 7723 66396
rect 7779 66394 7785 66396
rect 7539 66342 7541 66394
rect 7721 66342 7723 66394
rect 7477 66340 7483 66342
rect 7539 66340 7563 66342
rect 7619 66340 7643 66342
rect 7699 66340 7723 66342
rect 7779 66340 7785 66342
rect 7477 66320 7785 66340
rect 7477 65308 7785 65328
rect 7477 65306 7483 65308
rect 7539 65306 7563 65308
rect 7619 65306 7643 65308
rect 7699 65306 7723 65308
rect 7779 65306 7785 65308
rect 7539 65254 7541 65306
rect 7721 65254 7723 65306
rect 7477 65252 7483 65254
rect 7539 65252 7563 65254
rect 7619 65252 7643 65254
rect 7699 65252 7723 65254
rect 7779 65252 7785 65254
rect 7477 65232 7785 65252
rect 7477 64220 7785 64240
rect 7477 64218 7483 64220
rect 7539 64218 7563 64220
rect 7619 64218 7643 64220
rect 7699 64218 7723 64220
rect 7779 64218 7785 64220
rect 7539 64166 7541 64218
rect 7721 64166 7723 64218
rect 7477 64164 7483 64166
rect 7539 64164 7563 64166
rect 7619 64164 7643 64166
rect 7699 64164 7723 64166
rect 7779 64164 7785 64166
rect 7477 64144 7785 64164
rect 7477 63132 7785 63152
rect 7477 63130 7483 63132
rect 7539 63130 7563 63132
rect 7619 63130 7643 63132
rect 7699 63130 7723 63132
rect 7779 63130 7785 63132
rect 7539 63078 7541 63130
rect 7721 63078 7723 63130
rect 7477 63076 7483 63078
rect 7539 63076 7563 63078
rect 7619 63076 7643 63078
rect 7699 63076 7723 63078
rect 7779 63076 7785 63078
rect 7477 63056 7785 63076
rect 7477 62044 7785 62064
rect 7477 62042 7483 62044
rect 7539 62042 7563 62044
rect 7619 62042 7643 62044
rect 7699 62042 7723 62044
rect 7779 62042 7785 62044
rect 7539 61990 7541 62042
rect 7721 61990 7723 62042
rect 7477 61988 7483 61990
rect 7539 61988 7563 61990
rect 7619 61988 7643 61990
rect 7699 61988 7723 61990
rect 7779 61988 7785 61990
rect 7477 61968 7785 61988
rect 7477 60956 7785 60976
rect 7477 60954 7483 60956
rect 7539 60954 7563 60956
rect 7619 60954 7643 60956
rect 7699 60954 7723 60956
rect 7779 60954 7785 60956
rect 7539 60902 7541 60954
rect 7721 60902 7723 60954
rect 7477 60900 7483 60902
rect 7539 60900 7563 60902
rect 7619 60900 7643 60902
rect 7699 60900 7723 60902
rect 7779 60900 7785 60902
rect 7477 60880 7785 60900
rect 7477 59868 7785 59888
rect 7477 59866 7483 59868
rect 7539 59866 7563 59868
rect 7619 59866 7643 59868
rect 7699 59866 7723 59868
rect 7779 59866 7785 59868
rect 7539 59814 7541 59866
rect 7721 59814 7723 59866
rect 7477 59812 7483 59814
rect 7539 59812 7563 59814
rect 7619 59812 7643 59814
rect 7699 59812 7723 59814
rect 7779 59812 7785 59814
rect 7477 59792 7785 59812
rect 7477 58780 7785 58800
rect 7477 58778 7483 58780
rect 7539 58778 7563 58780
rect 7619 58778 7643 58780
rect 7699 58778 7723 58780
rect 7779 58778 7785 58780
rect 7539 58726 7541 58778
rect 7721 58726 7723 58778
rect 7477 58724 7483 58726
rect 7539 58724 7563 58726
rect 7619 58724 7643 58726
rect 7699 58724 7723 58726
rect 7779 58724 7785 58726
rect 7477 58704 7785 58724
rect 7477 57692 7785 57712
rect 7477 57690 7483 57692
rect 7539 57690 7563 57692
rect 7619 57690 7643 57692
rect 7699 57690 7723 57692
rect 7779 57690 7785 57692
rect 7539 57638 7541 57690
rect 7721 57638 7723 57690
rect 7477 57636 7483 57638
rect 7539 57636 7563 57638
rect 7619 57636 7643 57638
rect 7699 57636 7723 57638
rect 7779 57636 7785 57638
rect 7477 57616 7785 57636
rect 7196 57588 7248 57594
rect 7196 57530 7248 57536
rect 7024 46294 7144 46322
rect 7024 38758 7052 46294
rect 7208 45948 7236 57530
rect 7477 56604 7785 56624
rect 7477 56602 7483 56604
rect 7539 56602 7563 56604
rect 7619 56602 7643 56604
rect 7699 56602 7723 56604
rect 7779 56602 7785 56604
rect 7539 56550 7541 56602
rect 7721 56550 7723 56602
rect 7477 56548 7483 56550
rect 7539 56548 7563 56550
rect 7619 56548 7643 56550
rect 7699 56548 7723 56550
rect 7779 56548 7785 56550
rect 7477 56528 7785 56548
rect 7932 55820 7984 55826
rect 7932 55762 7984 55768
rect 7477 55516 7785 55536
rect 7477 55514 7483 55516
rect 7539 55514 7563 55516
rect 7619 55514 7643 55516
rect 7699 55514 7723 55516
rect 7779 55514 7785 55516
rect 7539 55462 7541 55514
rect 7721 55462 7723 55514
rect 7477 55460 7483 55462
rect 7539 55460 7563 55462
rect 7619 55460 7643 55462
rect 7699 55460 7723 55462
rect 7779 55460 7785 55462
rect 7477 55440 7785 55460
rect 7288 54596 7340 54602
rect 7288 54538 7340 54544
rect 7300 46102 7328 54538
rect 7477 54428 7785 54448
rect 7477 54426 7483 54428
rect 7539 54426 7563 54428
rect 7619 54426 7643 54428
rect 7699 54426 7723 54428
rect 7779 54426 7785 54428
rect 7539 54374 7541 54426
rect 7721 54374 7723 54426
rect 7477 54372 7483 54374
rect 7539 54372 7563 54374
rect 7619 54372 7643 54374
rect 7699 54372 7723 54374
rect 7779 54372 7785 54374
rect 7477 54352 7785 54372
rect 7477 53340 7785 53360
rect 7477 53338 7483 53340
rect 7539 53338 7563 53340
rect 7619 53338 7643 53340
rect 7699 53338 7723 53340
rect 7779 53338 7785 53340
rect 7539 53286 7541 53338
rect 7721 53286 7723 53338
rect 7477 53284 7483 53286
rect 7539 53284 7563 53286
rect 7619 53284 7643 53286
rect 7699 53284 7723 53286
rect 7779 53284 7785 53286
rect 7477 53264 7785 53284
rect 7380 52352 7432 52358
rect 7380 52294 7432 52300
rect 7392 46560 7420 52294
rect 7477 52252 7785 52272
rect 7477 52250 7483 52252
rect 7539 52250 7563 52252
rect 7619 52250 7643 52252
rect 7699 52250 7723 52252
rect 7779 52250 7785 52252
rect 7539 52198 7541 52250
rect 7721 52198 7723 52250
rect 7477 52196 7483 52198
rect 7539 52196 7563 52198
rect 7619 52196 7643 52198
rect 7699 52196 7723 52198
rect 7779 52196 7785 52198
rect 7477 52176 7785 52196
rect 7477 51164 7785 51184
rect 7477 51162 7483 51164
rect 7539 51162 7563 51164
rect 7619 51162 7643 51164
rect 7699 51162 7723 51164
rect 7779 51162 7785 51164
rect 7539 51110 7541 51162
rect 7721 51110 7723 51162
rect 7477 51108 7483 51110
rect 7539 51108 7563 51110
rect 7619 51108 7643 51110
rect 7699 51108 7723 51110
rect 7779 51108 7785 51110
rect 7477 51088 7785 51108
rect 7944 51074 7972 55762
rect 8024 53576 8076 53582
rect 8024 53518 8076 53524
rect 7852 51046 7972 51074
rect 7477 50076 7785 50096
rect 7477 50074 7483 50076
rect 7539 50074 7563 50076
rect 7619 50074 7643 50076
rect 7699 50074 7723 50076
rect 7779 50074 7785 50076
rect 7539 50022 7541 50074
rect 7721 50022 7723 50074
rect 7477 50020 7483 50022
rect 7539 50020 7563 50022
rect 7619 50020 7643 50022
rect 7699 50020 7723 50022
rect 7779 50020 7785 50022
rect 7477 50000 7785 50020
rect 7477 48988 7785 49008
rect 7477 48986 7483 48988
rect 7539 48986 7563 48988
rect 7619 48986 7643 48988
rect 7699 48986 7723 48988
rect 7779 48986 7785 48988
rect 7539 48934 7541 48986
rect 7721 48934 7723 48986
rect 7477 48932 7483 48934
rect 7539 48932 7563 48934
rect 7619 48932 7643 48934
rect 7699 48932 7723 48934
rect 7779 48932 7785 48934
rect 7477 48912 7785 48932
rect 7477 47900 7785 47920
rect 7477 47898 7483 47900
rect 7539 47898 7563 47900
rect 7619 47898 7643 47900
rect 7699 47898 7723 47900
rect 7779 47898 7785 47900
rect 7539 47846 7541 47898
rect 7721 47846 7723 47898
rect 7477 47844 7483 47846
rect 7539 47844 7563 47846
rect 7619 47844 7643 47846
rect 7699 47844 7723 47846
rect 7779 47844 7785 47846
rect 7477 47824 7785 47844
rect 7477 46812 7785 46832
rect 7477 46810 7483 46812
rect 7539 46810 7563 46812
rect 7619 46810 7643 46812
rect 7699 46810 7723 46812
rect 7779 46810 7785 46812
rect 7539 46758 7541 46810
rect 7721 46758 7723 46810
rect 7477 46756 7483 46758
rect 7539 46756 7563 46758
rect 7619 46756 7643 46758
rect 7699 46756 7723 46758
rect 7779 46756 7785 46758
rect 7477 46736 7785 46756
rect 7392 46532 7604 46560
rect 7288 46096 7340 46102
rect 7288 46038 7340 46044
rect 7380 46096 7432 46102
rect 7380 46038 7432 46044
rect 7576 46050 7604 46532
rect 7852 46170 7880 51046
rect 7932 47592 7984 47598
rect 7932 47534 7984 47540
rect 7944 46481 7972 47534
rect 7930 46472 7986 46481
rect 7930 46407 7986 46416
rect 8036 46322 8064 53518
rect 8116 53100 8168 53106
rect 8116 53042 8168 53048
rect 7944 46294 8064 46322
rect 7840 46164 7892 46170
rect 7840 46106 7892 46112
rect 7944 46102 7972 46294
rect 8128 46186 8156 53042
rect 8208 51808 8260 51814
rect 8208 51750 8260 51756
rect 8036 46158 8156 46186
rect 7932 46096 7984 46102
rect 7208 45920 7328 45948
rect 7104 45824 7156 45830
rect 7104 45766 7156 45772
rect 7196 45824 7248 45830
rect 7196 45766 7248 45772
rect 7012 38752 7064 38758
rect 7012 38694 7064 38700
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 7116 33522 7144 45766
rect 7104 33516 7156 33522
rect 7104 33458 7156 33464
rect 7208 31822 7236 45766
rect 7300 37738 7328 45920
rect 7288 37732 7340 37738
rect 7288 37674 7340 37680
rect 7196 31816 7248 31822
rect 7196 31758 7248 31764
rect 7392 27538 7420 46038
rect 7576 46022 7880 46050
rect 7932 46038 7984 46044
rect 7477 45724 7785 45744
rect 7477 45722 7483 45724
rect 7539 45722 7563 45724
rect 7619 45722 7643 45724
rect 7699 45722 7723 45724
rect 7779 45722 7785 45724
rect 7539 45670 7541 45722
rect 7721 45670 7723 45722
rect 7477 45668 7483 45670
rect 7539 45668 7563 45670
rect 7619 45668 7643 45670
rect 7699 45668 7723 45670
rect 7779 45668 7785 45670
rect 7477 45648 7785 45668
rect 7477 44636 7785 44656
rect 7477 44634 7483 44636
rect 7539 44634 7563 44636
rect 7619 44634 7643 44636
rect 7699 44634 7723 44636
rect 7779 44634 7785 44636
rect 7539 44582 7541 44634
rect 7721 44582 7723 44634
rect 7477 44580 7483 44582
rect 7539 44580 7563 44582
rect 7619 44580 7643 44582
rect 7699 44580 7723 44582
rect 7779 44580 7785 44582
rect 7477 44560 7785 44580
rect 7477 43548 7785 43568
rect 7477 43546 7483 43548
rect 7539 43546 7563 43548
rect 7619 43546 7643 43548
rect 7699 43546 7723 43548
rect 7779 43546 7785 43548
rect 7539 43494 7541 43546
rect 7721 43494 7723 43546
rect 7477 43492 7483 43494
rect 7539 43492 7563 43494
rect 7619 43492 7643 43494
rect 7699 43492 7723 43494
rect 7779 43492 7785 43494
rect 7477 43472 7785 43492
rect 7477 42460 7785 42480
rect 7477 42458 7483 42460
rect 7539 42458 7563 42460
rect 7619 42458 7643 42460
rect 7699 42458 7723 42460
rect 7779 42458 7785 42460
rect 7539 42406 7541 42458
rect 7721 42406 7723 42458
rect 7477 42404 7483 42406
rect 7539 42404 7563 42406
rect 7619 42404 7643 42406
rect 7699 42404 7723 42406
rect 7779 42404 7785 42406
rect 7477 42384 7785 42404
rect 7477 41372 7785 41392
rect 7477 41370 7483 41372
rect 7539 41370 7563 41372
rect 7619 41370 7643 41372
rect 7699 41370 7723 41372
rect 7779 41370 7785 41372
rect 7539 41318 7541 41370
rect 7721 41318 7723 41370
rect 7477 41316 7483 41318
rect 7539 41316 7563 41318
rect 7619 41316 7643 41318
rect 7699 41316 7723 41318
rect 7779 41316 7785 41318
rect 7477 41296 7785 41316
rect 7477 40284 7785 40304
rect 7477 40282 7483 40284
rect 7539 40282 7563 40284
rect 7619 40282 7643 40284
rect 7699 40282 7723 40284
rect 7779 40282 7785 40284
rect 7539 40230 7541 40282
rect 7721 40230 7723 40282
rect 7477 40228 7483 40230
rect 7539 40228 7563 40230
rect 7619 40228 7643 40230
rect 7699 40228 7723 40230
rect 7779 40228 7785 40230
rect 7477 40208 7785 40228
rect 7477 39196 7785 39216
rect 7477 39194 7483 39196
rect 7539 39194 7563 39196
rect 7619 39194 7643 39196
rect 7699 39194 7723 39196
rect 7779 39194 7785 39196
rect 7539 39142 7541 39194
rect 7721 39142 7723 39194
rect 7477 39140 7483 39142
rect 7539 39140 7563 39142
rect 7619 39140 7643 39142
rect 7699 39140 7723 39142
rect 7779 39140 7785 39142
rect 7477 39120 7785 39140
rect 7477 38108 7785 38128
rect 7477 38106 7483 38108
rect 7539 38106 7563 38108
rect 7619 38106 7643 38108
rect 7699 38106 7723 38108
rect 7779 38106 7785 38108
rect 7539 38054 7541 38106
rect 7721 38054 7723 38106
rect 7477 38052 7483 38054
rect 7539 38052 7563 38054
rect 7619 38052 7643 38054
rect 7699 38052 7723 38054
rect 7779 38052 7785 38054
rect 7477 38032 7785 38052
rect 7477 37020 7785 37040
rect 7477 37018 7483 37020
rect 7539 37018 7563 37020
rect 7619 37018 7643 37020
rect 7699 37018 7723 37020
rect 7779 37018 7785 37020
rect 7539 36966 7541 37018
rect 7721 36966 7723 37018
rect 7477 36964 7483 36966
rect 7539 36964 7563 36966
rect 7619 36964 7643 36966
rect 7699 36964 7723 36966
rect 7779 36964 7785 36966
rect 7477 36944 7785 36964
rect 7477 35932 7785 35952
rect 7477 35930 7483 35932
rect 7539 35930 7563 35932
rect 7619 35930 7643 35932
rect 7699 35930 7723 35932
rect 7779 35930 7785 35932
rect 7539 35878 7541 35930
rect 7721 35878 7723 35930
rect 7477 35876 7483 35878
rect 7539 35876 7563 35878
rect 7619 35876 7643 35878
rect 7699 35876 7723 35878
rect 7779 35876 7785 35878
rect 7477 35856 7785 35876
rect 7477 34844 7785 34864
rect 7477 34842 7483 34844
rect 7539 34842 7563 34844
rect 7619 34842 7643 34844
rect 7699 34842 7723 34844
rect 7779 34842 7785 34844
rect 7539 34790 7541 34842
rect 7721 34790 7723 34842
rect 7477 34788 7483 34790
rect 7539 34788 7563 34790
rect 7619 34788 7643 34790
rect 7699 34788 7723 34790
rect 7779 34788 7785 34790
rect 7477 34768 7785 34788
rect 7477 33756 7785 33776
rect 7477 33754 7483 33756
rect 7539 33754 7563 33756
rect 7619 33754 7643 33756
rect 7699 33754 7723 33756
rect 7779 33754 7785 33756
rect 7539 33702 7541 33754
rect 7721 33702 7723 33754
rect 7477 33700 7483 33702
rect 7539 33700 7563 33702
rect 7619 33700 7643 33702
rect 7699 33700 7723 33702
rect 7779 33700 7785 33702
rect 7477 33680 7785 33700
rect 7477 32668 7785 32688
rect 7477 32666 7483 32668
rect 7539 32666 7563 32668
rect 7619 32666 7643 32668
rect 7699 32666 7723 32668
rect 7779 32666 7785 32668
rect 7539 32614 7541 32666
rect 7721 32614 7723 32666
rect 7477 32612 7483 32614
rect 7539 32612 7563 32614
rect 7619 32612 7643 32614
rect 7699 32612 7723 32614
rect 7779 32612 7785 32614
rect 7477 32592 7785 32612
rect 7477 31580 7785 31600
rect 7477 31578 7483 31580
rect 7539 31578 7563 31580
rect 7619 31578 7643 31580
rect 7699 31578 7723 31580
rect 7779 31578 7785 31580
rect 7539 31526 7541 31578
rect 7721 31526 7723 31578
rect 7477 31524 7483 31526
rect 7539 31524 7563 31526
rect 7619 31524 7643 31526
rect 7699 31524 7723 31526
rect 7779 31524 7785 31526
rect 7477 31504 7785 31524
rect 7477 30492 7785 30512
rect 7477 30490 7483 30492
rect 7539 30490 7563 30492
rect 7619 30490 7643 30492
rect 7699 30490 7723 30492
rect 7779 30490 7785 30492
rect 7539 30438 7541 30490
rect 7721 30438 7723 30490
rect 7477 30436 7483 30438
rect 7539 30436 7563 30438
rect 7619 30436 7643 30438
rect 7699 30436 7723 30438
rect 7779 30436 7785 30438
rect 7477 30416 7785 30436
rect 7477 29404 7785 29424
rect 7477 29402 7483 29404
rect 7539 29402 7563 29404
rect 7619 29402 7643 29404
rect 7699 29402 7723 29404
rect 7779 29402 7785 29404
rect 7539 29350 7541 29402
rect 7721 29350 7723 29402
rect 7477 29348 7483 29350
rect 7539 29348 7563 29350
rect 7619 29348 7643 29350
rect 7699 29348 7723 29350
rect 7779 29348 7785 29350
rect 7477 29328 7785 29348
rect 7477 28316 7785 28336
rect 7477 28314 7483 28316
rect 7539 28314 7563 28316
rect 7619 28314 7643 28316
rect 7699 28314 7723 28316
rect 7779 28314 7785 28316
rect 7539 28262 7541 28314
rect 7721 28262 7723 28314
rect 7477 28260 7483 28262
rect 7539 28260 7563 28262
rect 7619 28260 7643 28262
rect 7699 28260 7723 28262
rect 7779 28260 7785 28262
rect 7477 28240 7785 28260
rect 7380 27532 7432 27538
rect 7380 27474 7432 27480
rect 7477 27228 7785 27248
rect 7477 27226 7483 27228
rect 7539 27226 7563 27228
rect 7619 27226 7643 27228
rect 7699 27226 7723 27228
rect 7779 27226 7785 27228
rect 7539 27174 7541 27226
rect 7721 27174 7723 27226
rect 7477 27172 7483 27174
rect 7539 27172 7563 27174
rect 7619 27172 7643 27174
rect 7699 27172 7723 27174
rect 7779 27172 7785 27174
rect 7477 27152 7785 27172
rect 7477 26140 7785 26160
rect 7477 26138 7483 26140
rect 7539 26138 7563 26140
rect 7619 26138 7643 26140
rect 7699 26138 7723 26140
rect 7779 26138 7785 26140
rect 7539 26086 7541 26138
rect 7721 26086 7723 26138
rect 7477 26084 7483 26086
rect 7539 26084 7563 26086
rect 7619 26084 7643 26086
rect 7699 26084 7723 26086
rect 7779 26084 7785 26086
rect 7477 26064 7785 26084
rect 7477 25052 7785 25072
rect 7477 25050 7483 25052
rect 7539 25050 7563 25052
rect 7619 25050 7643 25052
rect 7699 25050 7723 25052
rect 7779 25050 7785 25052
rect 7539 24998 7541 25050
rect 7721 24998 7723 25050
rect 7477 24996 7483 24998
rect 7539 24996 7563 24998
rect 7619 24996 7643 24998
rect 7699 24996 7723 24998
rect 7779 24996 7785 24998
rect 7477 24976 7785 24996
rect 7477 23964 7785 23984
rect 7477 23962 7483 23964
rect 7539 23962 7563 23964
rect 7619 23962 7643 23964
rect 7699 23962 7723 23964
rect 7779 23962 7785 23964
rect 7539 23910 7541 23962
rect 7721 23910 7723 23962
rect 7477 23908 7483 23910
rect 7539 23908 7563 23910
rect 7619 23908 7643 23910
rect 7699 23908 7723 23910
rect 7779 23908 7785 23910
rect 7477 23888 7785 23908
rect 7477 22876 7785 22896
rect 7477 22874 7483 22876
rect 7539 22874 7563 22876
rect 7619 22874 7643 22876
rect 7699 22874 7723 22876
rect 7779 22874 7785 22876
rect 7539 22822 7541 22874
rect 7721 22822 7723 22874
rect 7477 22820 7483 22822
rect 7539 22820 7563 22822
rect 7619 22820 7643 22822
rect 7699 22820 7723 22822
rect 7779 22820 7785 22822
rect 7477 22800 7785 22820
rect 7477 21788 7785 21808
rect 7477 21786 7483 21788
rect 7539 21786 7563 21788
rect 7619 21786 7643 21788
rect 7699 21786 7723 21788
rect 7779 21786 7785 21788
rect 7539 21734 7541 21786
rect 7721 21734 7723 21786
rect 7477 21732 7483 21734
rect 7539 21732 7563 21734
rect 7619 21732 7643 21734
rect 7699 21732 7723 21734
rect 7779 21732 7785 21734
rect 7477 21712 7785 21732
rect 7477 20700 7785 20720
rect 7477 20698 7483 20700
rect 7539 20698 7563 20700
rect 7619 20698 7643 20700
rect 7699 20698 7723 20700
rect 7779 20698 7785 20700
rect 7539 20646 7541 20698
rect 7721 20646 7723 20698
rect 7477 20644 7483 20646
rect 7539 20644 7563 20646
rect 7619 20644 7643 20646
rect 7699 20644 7723 20646
rect 7779 20644 7785 20646
rect 7477 20624 7785 20644
rect 7477 19612 7785 19632
rect 7477 19610 7483 19612
rect 7539 19610 7563 19612
rect 7619 19610 7643 19612
rect 7699 19610 7723 19612
rect 7779 19610 7785 19612
rect 7539 19558 7541 19610
rect 7721 19558 7723 19610
rect 7477 19556 7483 19558
rect 7539 19556 7563 19558
rect 7619 19556 7643 19558
rect 7699 19556 7723 19558
rect 7779 19556 7785 19558
rect 7477 19536 7785 19556
rect 7477 18524 7785 18544
rect 7477 18522 7483 18524
rect 7539 18522 7563 18524
rect 7619 18522 7643 18524
rect 7699 18522 7723 18524
rect 7779 18522 7785 18524
rect 7539 18470 7541 18522
rect 7721 18470 7723 18522
rect 7477 18468 7483 18470
rect 7539 18468 7563 18470
rect 7619 18468 7643 18470
rect 7699 18468 7723 18470
rect 7779 18468 7785 18470
rect 7477 18448 7785 18468
rect 7477 17436 7785 17456
rect 7477 17434 7483 17436
rect 7539 17434 7563 17436
rect 7619 17434 7643 17436
rect 7699 17434 7723 17436
rect 7779 17434 7785 17436
rect 7539 17382 7541 17434
rect 7721 17382 7723 17434
rect 7477 17380 7483 17382
rect 7539 17380 7563 17382
rect 7619 17380 7643 17382
rect 7699 17380 7723 17382
rect 7779 17380 7785 17382
rect 7477 17360 7785 17380
rect 7477 16348 7785 16368
rect 7477 16346 7483 16348
rect 7539 16346 7563 16348
rect 7619 16346 7643 16348
rect 7699 16346 7723 16348
rect 7779 16346 7785 16348
rect 7539 16294 7541 16346
rect 7721 16294 7723 16346
rect 7477 16292 7483 16294
rect 7539 16292 7563 16294
rect 7619 16292 7643 16294
rect 7699 16292 7723 16294
rect 7779 16292 7785 16294
rect 7477 16272 7785 16292
rect 7477 15260 7785 15280
rect 7477 15258 7483 15260
rect 7539 15258 7563 15260
rect 7619 15258 7643 15260
rect 7699 15258 7723 15260
rect 7779 15258 7785 15260
rect 7539 15206 7541 15258
rect 7721 15206 7723 15258
rect 7477 15204 7483 15206
rect 7539 15204 7563 15206
rect 7619 15204 7643 15206
rect 7699 15204 7723 15206
rect 7779 15204 7785 15206
rect 7477 15184 7785 15204
rect 7477 14172 7785 14192
rect 7477 14170 7483 14172
rect 7539 14170 7563 14172
rect 7619 14170 7643 14172
rect 7699 14170 7723 14172
rect 7779 14170 7785 14172
rect 7539 14118 7541 14170
rect 7721 14118 7723 14170
rect 7477 14116 7483 14118
rect 7539 14116 7563 14118
rect 7619 14116 7643 14118
rect 7699 14116 7723 14118
rect 7779 14116 7785 14118
rect 7477 14096 7785 14116
rect 7477 13084 7785 13104
rect 7477 13082 7483 13084
rect 7539 13082 7563 13084
rect 7619 13082 7643 13084
rect 7699 13082 7723 13084
rect 7779 13082 7785 13084
rect 7539 13030 7541 13082
rect 7721 13030 7723 13082
rect 7477 13028 7483 13030
rect 7539 13028 7563 13030
rect 7619 13028 7643 13030
rect 7699 13028 7723 13030
rect 7779 13028 7785 13030
rect 7477 13008 7785 13028
rect 7852 12442 7880 46022
rect 7932 45484 7984 45490
rect 7932 45426 7984 45432
rect 7944 36689 7972 45426
rect 7930 36680 7986 36689
rect 7930 36615 7986 36624
rect 7932 36576 7984 36582
rect 7932 36518 7984 36524
rect 7944 15094 7972 36518
rect 8036 29102 8064 46158
rect 8114 46064 8170 46073
rect 8114 45999 8170 46008
rect 8128 36582 8156 45999
rect 8116 36576 8168 36582
rect 8116 36518 8168 36524
rect 8114 36408 8170 36417
rect 8114 36343 8170 36352
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7477 11996 7785 12016
rect 7477 11994 7483 11996
rect 7539 11994 7563 11996
rect 7619 11994 7643 11996
rect 7699 11994 7723 11996
rect 7779 11994 7785 11996
rect 7539 11942 7541 11994
rect 7721 11942 7723 11994
rect 7477 11940 7483 11942
rect 7539 11940 7563 11942
rect 7619 11940 7643 11942
rect 7699 11940 7723 11942
rect 7779 11940 7785 11942
rect 7477 11920 7785 11940
rect 7477 10908 7785 10928
rect 7477 10906 7483 10908
rect 7539 10906 7563 10908
rect 7619 10906 7643 10908
rect 7699 10906 7723 10908
rect 7779 10906 7785 10908
rect 7539 10854 7541 10906
rect 7721 10854 7723 10906
rect 7477 10852 7483 10854
rect 7539 10852 7563 10854
rect 7619 10852 7643 10854
rect 7699 10852 7723 10854
rect 7779 10852 7785 10854
rect 7477 10832 7785 10852
rect 7477 9820 7785 9840
rect 7477 9818 7483 9820
rect 7539 9818 7563 9820
rect 7619 9818 7643 9820
rect 7699 9818 7723 9820
rect 7779 9818 7785 9820
rect 7539 9766 7541 9818
rect 7721 9766 7723 9818
rect 7477 9764 7483 9766
rect 7539 9764 7563 9766
rect 7619 9764 7643 9766
rect 7699 9764 7723 9766
rect 7779 9764 7785 9766
rect 7477 9744 7785 9764
rect 7477 8732 7785 8752
rect 7477 8730 7483 8732
rect 7539 8730 7563 8732
rect 7619 8730 7643 8732
rect 7699 8730 7723 8732
rect 7779 8730 7785 8732
rect 7539 8678 7541 8730
rect 7721 8678 7723 8730
rect 7477 8676 7483 8678
rect 7539 8676 7563 8678
rect 7619 8676 7643 8678
rect 7699 8676 7723 8678
rect 7779 8676 7785 8678
rect 7477 8656 7785 8676
rect 7477 7644 7785 7664
rect 7477 7642 7483 7644
rect 7539 7642 7563 7644
rect 7619 7642 7643 7644
rect 7699 7642 7723 7644
rect 7779 7642 7785 7644
rect 7539 7590 7541 7642
rect 7721 7590 7723 7642
rect 7477 7588 7483 7590
rect 7539 7588 7563 7590
rect 7619 7588 7643 7590
rect 7699 7588 7723 7590
rect 7779 7588 7785 7590
rect 7477 7568 7785 7588
rect 7477 6556 7785 6576
rect 7477 6554 7483 6556
rect 7539 6554 7563 6556
rect 7619 6554 7643 6556
rect 7699 6554 7723 6556
rect 7779 6554 7785 6556
rect 7539 6502 7541 6554
rect 7721 6502 7723 6554
rect 7477 6500 7483 6502
rect 7539 6500 7563 6502
rect 7619 6500 7643 6502
rect 7699 6500 7723 6502
rect 7779 6500 7785 6502
rect 7477 6480 7785 6500
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 7477 5468 7785 5488
rect 7477 5466 7483 5468
rect 7539 5466 7563 5468
rect 7619 5466 7643 5468
rect 7699 5466 7723 5468
rect 7779 5466 7785 5468
rect 7539 5414 7541 5466
rect 7721 5414 7723 5466
rect 7477 5412 7483 5414
rect 7539 5412 7563 5414
rect 7619 5412 7643 5414
rect 7699 5412 7723 5414
rect 7779 5412 7785 5414
rect 7477 5392 7785 5412
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5845 3836 6153 3856
rect 5845 3834 5851 3836
rect 5907 3834 5931 3836
rect 5987 3834 6011 3836
rect 6067 3834 6091 3836
rect 6147 3834 6153 3836
rect 5907 3782 5909 3834
rect 6089 3782 6091 3834
rect 5845 3780 5851 3782
rect 5907 3780 5931 3782
rect 5987 3780 6011 3782
rect 6067 3780 6091 3782
rect 6147 3780 6153 3782
rect 5845 3760 6153 3780
rect 4213 3292 4521 3312
rect 4213 3290 4219 3292
rect 4275 3290 4299 3292
rect 4355 3290 4379 3292
rect 4435 3290 4459 3292
rect 4515 3290 4521 3292
rect 4275 3238 4277 3290
rect 4457 3238 4459 3290
rect 4213 3236 4219 3238
rect 4275 3236 4299 3238
rect 4355 3236 4379 3238
rect 4435 3236 4459 3238
rect 4515 3236 4521 3238
rect 4213 3216 4521 3236
rect 6380 3058 6408 4966
rect 7477 4380 7785 4400
rect 7477 4378 7483 4380
rect 7539 4378 7563 4380
rect 7619 4378 7643 4380
rect 7699 4378 7723 4380
rect 7779 4378 7785 4380
rect 7539 4326 7541 4378
rect 7721 4326 7723 4378
rect 7477 4324 7483 4326
rect 7539 4324 7563 4326
rect 7619 4324 7643 4326
rect 7699 4324 7723 4326
rect 7779 4324 7785 4326
rect 7477 4304 7785 4324
rect 8128 3670 8156 36343
rect 8220 11354 8248 51750
rect 8312 43994 8340 74598
rect 9109 74556 9417 74576
rect 9109 74554 9115 74556
rect 9171 74554 9195 74556
rect 9251 74554 9275 74556
rect 9331 74554 9355 74556
rect 9411 74554 9417 74556
rect 9171 74502 9173 74554
rect 9353 74502 9355 74554
rect 9109 74500 9115 74502
rect 9171 74500 9195 74502
rect 9251 74500 9275 74502
rect 9331 74500 9355 74502
rect 9411 74500 9417 74502
rect 9109 74480 9417 74500
rect 10140 74248 10192 74254
rect 10138 74216 10140 74225
rect 10192 74216 10194 74225
rect 10138 74151 10194 74160
rect 9772 74112 9824 74118
rect 9772 74054 9824 74060
rect 9109 73468 9417 73488
rect 9109 73466 9115 73468
rect 9171 73466 9195 73468
rect 9251 73466 9275 73468
rect 9331 73466 9355 73468
rect 9411 73466 9417 73468
rect 9171 73414 9173 73466
rect 9353 73414 9355 73466
rect 9109 73412 9115 73414
rect 9171 73412 9195 73414
rect 9251 73412 9275 73414
rect 9331 73412 9355 73414
rect 9411 73412 9417 73414
rect 9109 73392 9417 73412
rect 9109 72380 9417 72400
rect 9109 72378 9115 72380
rect 9171 72378 9195 72380
rect 9251 72378 9275 72380
rect 9331 72378 9355 72380
rect 9411 72378 9417 72380
rect 9171 72326 9173 72378
rect 9353 72326 9355 72378
rect 9109 72324 9115 72326
rect 9171 72324 9195 72326
rect 9251 72324 9275 72326
rect 9331 72324 9355 72326
rect 9411 72324 9417 72326
rect 9109 72304 9417 72324
rect 9784 71738 9812 74054
rect 10140 73772 10192 73778
rect 10140 73714 10192 73720
rect 9956 73704 10008 73710
rect 9956 73646 10008 73652
rect 9968 72282 9996 73646
rect 10152 73409 10180 73714
rect 10138 73400 10194 73409
rect 10138 73335 10194 73344
rect 10140 73160 10192 73166
rect 10140 73102 10192 73108
rect 10152 72729 10180 73102
rect 10138 72720 10194 72729
rect 10138 72655 10194 72664
rect 9956 72276 10008 72282
rect 9956 72218 10008 72224
rect 10140 72072 10192 72078
rect 10140 72014 10192 72020
rect 9864 72004 9916 72010
rect 9864 71946 9916 71952
rect 9772 71732 9824 71738
rect 9772 71674 9824 71680
rect 9109 71292 9417 71312
rect 9109 71290 9115 71292
rect 9171 71290 9195 71292
rect 9251 71290 9275 71292
rect 9331 71290 9355 71292
rect 9411 71290 9417 71292
rect 9171 71238 9173 71290
rect 9353 71238 9355 71290
rect 9109 71236 9115 71238
rect 9171 71236 9195 71238
rect 9251 71236 9275 71238
rect 9331 71236 9355 71238
rect 9411 71236 9417 71238
rect 9109 71216 9417 71236
rect 9876 70650 9904 71946
rect 10152 71913 10180 72014
rect 10138 71904 10194 71913
rect 10138 71839 10194 71848
rect 10140 71596 10192 71602
rect 10140 71538 10192 71544
rect 10152 71097 10180 71538
rect 10138 71088 10194 71097
rect 10138 71023 10194 71032
rect 9864 70644 9916 70650
rect 9864 70586 9916 70592
rect 10140 70508 10192 70514
rect 10140 70450 10192 70456
rect 10152 70417 10180 70450
rect 10138 70408 10194 70417
rect 10138 70343 10194 70352
rect 9109 70204 9417 70224
rect 9109 70202 9115 70204
rect 9171 70202 9195 70204
rect 9251 70202 9275 70204
rect 9331 70202 9355 70204
rect 9411 70202 9417 70204
rect 9171 70150 9173 70202
rect 9353 70150 9355 70202
rect 9109 70148 9115 70150
rect 9171 70148 9195 70150
rect 9251 70148 9275 70150
rect 9331 70148 9355 70150
rect 9411 70148 9417 70150
rect 9109 70128 9417 70148
rect 10140 69896 10192 69902
rect 10140 69838 10192 69844
rect 9956 69760 10008 69766
rect 9956 69702 10008 69708
rect 9968 69494 9996 69702
rect 10152 69601 10180 69838
rect 10138 69592 10194 69601
rect 10138 69527 10194 69536
rect 9956 69488 10008 69494
rect 9956 69430 10008 69436
rect 10140 69420 10192 69426
rect 10140 69362 10192 69368
rect 9956 69216 10008 69222
rect 9956 69158 10008 69164
rect 9109 69116 9417 69136
rect 9109 69114 9115 69116
rect 9171 69114 9195 69116
rect 9251 69114 9275 69116
rect 9331 69114 9355 69116
rect 9411 69114 9417 69116
rect 9171 69062 9173 69114
rect 9353 69062 9355 69114
rect 9109 69060 9115 69062
rect 9171 69060 9195 69062
rect 9251 69060 9275 69062
rect 9331 69060 9355 69062
rect 9411 69060 9417 69062
rect 9109 69040 9417 69060
rect 9968 68406 9996 69158
rect 10152 68921 10180 69362
rect 10138 68912 10194 68921
rect 10138 68847 10194 68856
rect 9956 68400 10008 68406
rect 9956 68342 10008 68348
rect 10140 68332 10192 68338
rect 10140 68274 10192 68280
rect 8484 68128 8536 68134
rect 10152 68105 10180 68274
rect 8484 68070 8536 68076
rect 10138 68096 10194 68105
rect 8392 55276 8444 55282
rect 8392 55218 8444 55224
rect 8300 43988 8352 43994
rect 8300 43930 8352 43936
rect 8404 35222 8432 55218
rect 8496 39846 8524 68070
rect 9109 68028 9417 68048
rect 10138 68031 10194 68040
rect 9109 68026 9115 68028
rect 9171 68026 9195 68028
rect 9251 68026 9275 68028
rect 9331 68026 9355 68028
rect 9411 68026 9417 68028
rect 9171 67974 9173 68026
rect 9353 67974 9355 68026
rect 9109 67972 9115 67974
rect 9171 67972 9195 67974
rect 9251 67972 9275 67974
rect 9331 67972 9355 67974
rect 9411 67972 9417 67974
rect 9109 67952 9417 67972
rect 9956 67584 10008 67590
rect 9956 67526 10008 67532
rect 10140 67584 10192 67590
rect 10140 67526 10192 67532
rect 9968 67318 9996 67526
rect 9956 67312 10008 67318
rect 10152 67289 10180 67526
rect 9956 67254 10008 67260
rect 10138 67280 10194 67289
rect 10138 67215 10194 67224
rect 9109 66940 9417 66960
rect 9109 66938 9115 66940
rect 9171 66938 9195 66940
rect 9251 66938 9275 66940
rect 9331 66938 9355 66940
rect 9411 66938 9417 66940
rect 9171 66886 9173 66938
rect 9353 66886 9355 66938
rect 9109 66884 9115 66886
rect 9171 66884 9195 66886
rect 9251 66884 9275 66886
rect 9331 66884 9355 66886
rect 9411 66884 9417 66886
rect 9109 66864 9417 66884
rect 10140 66632 10192 66638
rect 10138 66600 10140 66609
rect 10192 66600 10194 66609
rect 10138 66535 10194 66544
rect 9956 66496 10008 66502
rect 9956 66438 10008 66444
rect 9864 65952 9916 65958
rect 9864 65894 9916 65900
rect 9109 65852 9417 65872
rect 9109 65850 9115 65852
rect 9171 65850 9195 65852
rect 9251 65850 9275 65852
rect 9331 65850 9355 65852
rect 9411 65850 9417 65852
rect 9171 65798 9173 65850
rect 9353 65798 9355 65850
rect 9109 65796 9115 65798
rect 9171 65796 9195 65798
rect 9251 65796 9275 65798
rect 9331 65796 9355 65798
rect 9411 65796 9417 65798
rect 9109 65776 9417 65796
rect 9772 65408 9824 65414
rect 9772 65350 9824 65356
rect 9109 64764 9417 64784
rect 9109 64762 9115 64764
rect 9171 64762 9195 64764
rect 9251 64762 9275 64764
rect 9331 64762 9355 64764
rect 9411 64762 9417 64764
rect 9171 64710 9173 64762
rect 9353 64710 9355 64762
rect 9109 64708 9115 64710
rect 9171 64708 9195 64710
rect 9251 64708 9275 64710
rect 9331 64708 9355 64710
rect 9411 64708 9417 64710
rect 9109 64688 9417 64708
rect 9109 63676 9417 63696
rect 9109 63674 9115 63676
rect 9171 63674 9195 63676
rect 9251 63674 9275 63676
rect 9331 63674 9355 63676
rect 9411 63674 9417 63676
rect 9171 63622 9173 63674
rect 9353 63622 9355 63674
rect 9109 63620 9115 63622
rect 9171 63620 9195 63622
rect 9251 63620 9275 63622
rect 9331 63620 9355 63622
rect 9411 63620 9417 63622
rect 9109 63600 9417 63620
rect 8576 63504 8628 63510
rect 8576 63446 8628 63452
rect 8484 39840 8536 39846
rect 8484 39782 8536 39788
rect 8588 36242 8616 63446
rect 9784 62966 9812 65350
rect 9876 64122 9904 65894
rect 9968 65142 9996 66438
rect 10140 66156 10192 66162
rect 10140 66098 10192 66104
rect 10152 65793 10180 66098
rect 10138 65784 10194 65793
rect 10138 65719 10194 65728
rect 10140 65544 10192 65550
rect 10140 65486 10192 65492
rect 9956 65136 10008 65142
rect 10152 65113 10180 65486
rect 9956 65078 10008 65084
rect 10138 65104 10194 65113
rect 10138 65039 10194 65048
rect 10140 64456 10192 64462
rect 10140 64398 10192 64404
rect 10152 64297 10180 64398
rect 10138 64288 10194 64297
rect 10138 64223 10194 64232
rect 9864 64116 9916 64122
rect 9864 64058 9916 64064
rect 10140 63912 10192 63918
rect 10140 63854 10192 63860
rect 10152 63481 10180 63854
rect 10138 63472 10194 63481
rect 10138 63407 10194 63416
rect 9956 63300 10008 63306
rect 9956 63242 10008 63248
rect 9968 63034 9996 63242
rect 9956 63028 10008 63034
rect 9956 62970 10008 62976
rect 9772 62960 9824 62966
rect 9772 62902 9824 62908
rect 10140 62892 10192 62898
rect 10140 62834 10192 62840
rect 10152 62801 10180 62834
rect 10138 62792 10194 62801
rect 10138 62727 10194 62736
rect 9109 62588 9417 62608
rect 9109 62586 9115 62588
rect 9171 62586 9195 62588
rect 9251 62586 9275 62588
rect 9331 62586 9355 62588
rect 9411 62586 9417 62588
rect 9171 62534 9173 62586
rect 9353 62534 9355 62586
rect 9109 62532 9115 62534
rect 9171 62532 9195 62534
rect 9251 62532 9275 62534
rect 9331 62532 9355 62534
rect 9411 62532 9417 62534
rect 9109 62512 9417 62532
rect 9680 62348 9732 62354
rect 9680 62290 9732 62296
rect 9109 61500 9417 61520
rect 9109 61498 9115 61500
rect 9171 61498 9195 61500
rect 9251 61498 9275 61500
rect 9331 61498 9355 61500
rect 9411 61498 9417 61500
rect 9171 61446 9173 61498
rect 9353 61446 9355 61498
rect 9109 61444 9115 61446
rect 9171 61444 9195 61446
rect 9251 61444 9275 61446
rect 9331 61444 9355 61446
rect 9411 61444 9417 61446
rect 9109 61424 9417 61444
rect 9109 60412 9417 60432
rect 9109 60410 9115 60412
rect 9171 60410 9195 60412
rect 9251 60410 9275 60412
rect 9331 60410 9355 60412
rect 9411 60410 9417 60412
rect 9171 60358 9173 60410
rect 9353 60358 9355 60410
rect 9109 60356 9115 60358
rect 9171 60356 9195 60358
rect 9251 60356 9275 60358
rect 9331 60356 9355 60358
rect 9411 60356 9417 60358
rect 9109 60336 9417 60356
rect 9692 60314 9720 62290
rect 10140 62280 10192 62286
rect 10140 62222 10192 62228
rect 10152 61985 10180 62222
rect 10138 61976 10194 61985
rect 10138 61911 10194 61920
rect 10140 61804 10192 61810
rect 10140 61746 10192 61752
rect 9772 61736 9824 61742
rect 9772 61678 9824 61684
rect 9784 60586 9812 61678
rect 9956 61600 10008 61606
rect 9956 61542 10008 61548
rect 9864 61124 9916 61130
rect 9864 61066 9916 61072
rect 9772 60580 9824 60586
rect 9772 60522 9824 60528
rect 9680 60308 9732 60314
rect 9680 60250 9732 60256
rect 9109 59324 9417 59344
rect 9109 59322 9115 59324
rect 9171 59322 9195 59324
rect 9251 59322 9275 59324
rect 9331 59322 9355 59324
rect 9411 59322 9417 59324
rect 9171 59270 9173 59322
rect 9353 59270 9355 59322
rect 9109 59268 9115 59270
rect 9171 59268 9195 59270
rect 9251 59268 9275 59270
rect 9331 59268 9355 59270
rect 9411 59268 9417 59270
rect 9109 59248 9417 59268
rect 9876 59226 9904 61066
rect 9968 60790 9996 61542
rect 10152 61305 10180 61746
rect 10138 61296 10194 61305
rect 10138 61231 10194 61240
rect 9956 60784 10008 60790
rect 9956 60726 10008 60732
rect 10140 60716 10192 60722
rect 10140 60658 10192 60664
rect 10152 60489 10180 60658
rect 10138 60480 10194 60489
rect 10138 60415 10194 60424
rect 10140 60104 10192 60110
rect 10140 60046 10192 60052
rect 10152 59673 10180 60046
rect 10138 59664 10194 59673
rect 10138 59599 10194 59608
rect 9864 59220 9916 59226
rect 9864 59162 9916 59168
rect 10140 59016 10192 59022
rect 10138 58984 10140 58993
rect 10192 58984 10194 58993
rect 10138 58919 10194 58928
rect 10140 58540 10192 58546
rect 10140 58482 10192 58488
rect 9956 58336 10008 58342
rect 9956 58278 10008 58284
rect 9109 58236 9417 58256
rect 9109 58234 9115 58236
rect 9171 58234 9195 58236
rect 9251 58234 9275 58236
rect 9331 58234 9355 58236
rect 9411 58234 9417 58236
rect 9171 58182 9173 58234
rect 9353 58182 9355 58234
rect 9109 58180 9115 58182
rect 9171 58180 9195 58182
rect 9251 58180 9275 58182
rect 9331 58180 9355 58182
rect 9411 58180 9417 58182
rect 9109 58160 9417 58180
rect 9968 57390 9996 58278
rect 10152 58177 10180 58482
rect 10138 58168 10194 58177
rect 10138 58103 10194 58112
rect 10140 57928 10192 57934
rect 10140 57870 10192 57876
rect 10152 57497 10180 57870
rect 10138 57488 10194 57497
rect 10138 57423 10194 57432
rect 9956 57384 10008 57390
rect 9956 57326 10008 57332
rect 9109 57148 9417 57168
rect 9109 57146 9115 57148
rect 9171 57146 9195 57148
rect 9251 57146 9275 57148
rect 9331 57146 9355 57148
rect 9411 57146 9417 57148
rect 9171 57094 9173 57146
rect 9353 57094 9355 57146
rect 9109 57092 9115 57094
rect 9171 57092 9195 57094
rect 9251 57092 9275 57094
rect 9331 57092 9355 57094
rect 9411 57092 9417 57094
rect 9109 57072 9417 57092
rect 10140 56840 10192 56846
rect 10140 56782 10192 56788
rect 8760 56704 8812 56710
rect 10152 56681 10180 56782
rect 8760 56646 8812 56652
rect 10138 56672 10194 56681
rect 8668 55752 8720 55758
rect 8668 55694 8720 55700
rect 8576 36236 8628 36242
rect 8576 36178 8628 36184
rect 8392 35216 8444 35222
rect 8392 35158 8444 35164
rect 8680 34678 8708 55694
rect 8772 37126 8800 56646
rect 10138 56607 10194 56616
rect 8852 56364 8904 56370
rect 8852 56306 8904 56312
rect 10140 56364 10192 56370
rect 10140 56306 10192 56312
rect 8760 37120 8812 37126
rect 8760 37062 8812 37068
rect 8864 35562 8892 56306
rect 9956 56160 10008 56166
rect 9956 56102 10008 56108
rect 9109 56060 9417 56080
rect 9109 56058 9115 56060
rect 9171 56058 9195 56060
rect 9251 56058 9275 56060
rect 9331 56058 9355 56060
rect 9411 56058 9417 56060
rect 9171 56006 9173 56058
rect 9353 56006 9355 56058
rect 9109 56004 9115 56006
rect 9171 56004 9195 56006
rect 9251 56004 9275 56006
rect 9331 56004 9355 56006
rect 9411 56004 9417 56006
rect 9109 55984 9417 56004
rect 9968 55418 9996 56102
rect 10152 55865 10180 56306
rect 10138 55856 10194 55865
rect 10138 55791 10194 55800
rect 9956 55412 10008 55418
rect 9956 55354 10008 55360
rect 10140 55276 10192 55282
rect 10140 55218 10192 55224
rect 10152 55185 10180 55218
rect 10138 55176 10194 55185
rect 10138 55111 10194 55120
rect 9956 55072 10008 55078
rect 9956 55014 10008 55020
rect 9109 54972 9417 54992
rect 9109 54970 9115 54972
rect 9171 54970 9195 54972
rect 9251 54970 9275 54972
rect 9331 54970 9355 54972
rect 9411 54970 9417 54972
rect 9171 54918 9173 54970
rect 9353 54918 9355 54970
rect 9109 54916 9115 54918
rect 9171 54916 9195 54918
rect 9251 54916 9275 54918
rect 9331 54916 9355 54918
rect 9411 54916 9417 54918
rect 9109 54896 9417 54916
rect 9772 54188 9824 54194
rect 9772 54130 9824 54136
rect 9109 53884 9417 53904
rect 9109 53882 9115 53884
rect 9171 53882 9195 53884
rect 9251 53882 9275 53884
rect 9331 53882 9355 53884
rect 9411 53882 9417 53884
rect 9171 53830 9173 53882
rect 9353 53830 9355 53882
rect 9109 53828 9115 53830
rect 9171 53828 9195 53830
rect 9251 53828 9275 53830
rect 9331 53828 9355 53830
rect 9411 53828 9417 53830
rect 9109 53808 9417 53828
rect 9109 52796 9417 52816
rect 9109 52794 9115 52796
rect 9171 52794 9195 52796
rect 9251 52794 9275 52796
rect 9331 52794 9355 52796
rect 9411 52794 9417 52796
rect 9171 52742 9173 52794
rect 9353 52742 9355 52794
rect 9109 52740 9115 52742
rect 9171 52740 9195 52742
rect 9251 52740 9275 52742
rect 9331 52740 9355 52742
rect 9411 52740 9417 52742
rect 9109 52720 9417 52740
rect 9784 52698 9812 54130
rect 9968 53514 9996 55014
rect 10140 54664 10192 54670
rect 10140 54606 10192 54612
rect 10152 54369 10180 54606
rect 10138 54360 10194 54369
rect 10138 54295 10194 54304
rect 10048 53984 10100 53990
rect 10048 53926 10100 53932
rect 10060 53689 10088 53926
rect 10046 53680 10102 53689
rect 10046 53615 10102 53624
rect 9956 53508 10008 53514
rect 9956 53450 10008 53456
rect 9864 53100 9916 53106
rect 9864 53042 9916 53048
rect 9772 52692 9824 52698
rect 9772 52634 9824 52640
rect 9876 52154 9904 53042
rect 10048 52896 10100 52902
rect 10046 52864 10048 52873
rect 10100 52864 10102 52873
rect 10046 52799 10102 52808
rect 10048 52352 10100 52358
rect 10048 52294 10100 52300
rect 9864 52148 9916 52154
rect 9864 52090 9916 52096
rect 10060 52057 10088 52294
rect 10046 52048 10102 52057
rect 10046 51983 10102 51992
rect 9109 51708 9417 51728
rect 9109 51706 9115 51708
rect 9171 51706 9195 51708
rect 9251 51706 9275 51708
rect 9331 51706 9355 51708
rect 9411 51706 9417 51708
rect 9171 51654 9173 51706
rect 9353 51654 9355 51706
rect 9109 51652 9115 51654
rect 9171 51652 9195 51654
rect 9251 51652 9275 51654
rect 9331 51652 9355 51654
rect 9411 51652 9417 51654
rect 9109 51632 9417 51652
rect 9864 51400 9916 51406
rect 9864 51342 9916 51348
rect 10046 51368 10102 51377
rect 9109 50620 9417 50640
rect 9109 50618 9115 50620
rect 9171 50618 9195 50620
rect 9251 50618 9275 50620
rect 9331 50618 9355 50620
rect 9411 50618 9417 50620
rect 9171 50566 9173 50618
rect 9353 50566 9355 50618
rect 9109 50564 9115 50566
rect 9171 50564 9195 50566
rect 9251 50564 9275 50566
rect 9331 50564 9355 50566
rect 9411 50564 9417 50566
rect 9109 50544 9417 50564
rect 9876 50522 9904 51342
rect 10046 51303 10102 51312
rect 10060 51270 10088 51303
rect 10048 51264 10100 51270
rect 10048 51206 10100 51212
rect 10048 50720 10100 50726
rect 10048 50662 10100 50668
rect 10060 50561 10088 50662
rect 10046 50552 10102 50561
rect 9864 50516 9916 50522
rect 10046 50487 10102 50496
rect 9864 50458 9916 50464
rect 10968 50380 11020 50386
rect 10968 50322 11020 50328
rect 10048 50176 10100 50182
rect 10048 50118 10100 50124
rect 10060 49881 10088 50118
rect 10046 49872 10102 49881
rect 10980 49842 11008 50322
rect 10046 49807 10102 49816
rect 10968 49836 11020 49842
rect 10968 49778 11020 49784
rect 9680 49768 9732 49774
rect 9680 49710 9732 49716
rect 9109 49532 9417 49552
rect 9109 49530 9115 49532
rect 9171 49530 9195 49532
rect 9251 49530 9275 49532
rect 9331 49530 9355 49532
rect 9411 49530 9417 49532
rect 9171 49478 9173 49530
rect 9353 49478 9355 49530
rect 9109 49476 9115 49478
rect 9171 49476 9195 49478
rect 9251 49476 9275 49478
rect 9331 49476 9355 49478
rect 9411 49476 9417 49478
rect 9109 49456 9417 49476
rect 9588 49224 9640 49230
rect 9588 49166 9640 49172
rect 9109 48444 9417 48464
rect 9109 48442 9115 48444
rect 9171 48442 9195 48444
rect 9251 48442 9275 48444
rect 9331 48442 9355 48444
rect 9411 48442 9417 48444
rect 9171 48390 9173 48442
rect 9353 48390 9355 48442
rect 9109 48388 9115 48390
rect 9171 48388 9195 48390
rect 9251 48388 9275 48390
rect 9331 48388 9355 48390
rect 9411 48388 9417 48390
rect 9109 48368 9417 48388
rect 9036 47524 9088 47530
rect 9036 47466 9088 47472
rect 8944 47116 8996 47122
rect 8944 47058 8996 47064
rect 8852 35556 8904 35562
rect 8852 35498 8904 35504
rect 8668 34672 8720 34678
rect 8668 34614 8720 34620
rect 8956 14278 8984 47058
rect 9048 15162 9076 47466
rect 9109 47356 9417 47376
rect 9109 47354 9115 47356
rect 9171 47354 9195 47356
rect 9251 47354 9275 47356
rect 9331 47354 9355 47356
rect 9411 47354 9417 47356
rect 9171 47302 9173 47354
rect 9353 47302 9355 47354
rect 9109 47300 9115 47302
rect 9171 47300 9195 47302
rect 9251 47300 9275 47302
rect 9331 47300 9355 47302
rect 9411 47300 9417 47302
rect 9109 47280 9417 47300
rect 9600 46714 9628 49166
rect 9692 47666 9720 49710
rect 9864 49088 9916 49094
rect 10048 49088 10100 49094
rect 9864 49030 9916 49036
rect 10046 49056 10048 49065
rect 10100 49056 10102 49065
rect 9772 48748 9824 48754
rect 9772 48690 9824 48696
rect 9784 48278 9812 48690
rect 9772 48272 9824 48278
rect 9772 48214 9824 48220
rect 9680 47660 9732 47666
rect 9680 47602 9732 47608
rect 9588 46708 9640 46714
rect 9588 46650 9640 46656
rect 9876 46578 9904 49030
rect 10046 48991 10102 49000
rect 10048 48544 10100 48550
rect 10048 48486 10100 48492
rect 10060 48249 10088 48486
rect 10046 48240 10102 48249
rect 10046 48175 10102 48184
rect 10046 47560 10102 47569
rect 10046 47495 10048 47504
rect 10100 47495 10102 47504
rect 10048 47466 10100 47472
rect 10048 46912 10100 46918
rect 10048 46854 10100 46860
rect 10060 46753 10088 46854
rect 10046 46744 10102 46753
rect 10046 46679 10102 46688
rect 9864 46572 9916 46578
rect 9864 46514 9916 46520
rect 10048 46368 10100 46374
rect 10048 46310 10100 46316
rect 9109 46268 9417 46288
rect 9109 46266 9115 46268
rect 9171 46266 9195 46268
rect 9251 46266 9275 46268
rect 9331 46266 9355 46268
rect 9411 46266 9417 46268
rect 9171 46214 9173 46266
rect 9353 46214 9355 46266
rect 9109 46212 9115 46214
rect 9171 46212 9195 46214
rect 9251 46212 9275 46214
rect 9331 46212 9355 46214
rect 9411 46212 9417 46214
rect 9109 46192 9417 46212
rect 10060 46073 10088 46310
rect 10046 46064 10102 46073
rect 10046 45999 10102 46008
rect 10048 45280 10100 45286
rect 10046 45248 10048 45257
rect 10100 45248 10102 45257
rect 9109 45180 9417 45200
rect 10046 45183 10102 45192
rect 9109 45178 9115 45180
rect 9171 45178 9195 45180
rect 9251 45178 9275 45180
rect 9331 45178 9355 45180
rect 9411 45178 9417 45180
rect 9171 45126 9173 45178
rect 9353 45126 9355 45178
rect 9109 45124 9115 45126
rect 9171 45124 9195 45126
rect 9251 45124 9275 45126
rect 9331 45124 9355 45126
rect 9411 45124 9417 45126
rect 9109 45104 9417 45124
rect 9864 44736 9916 44742
rect 9864 44678 9916 44684
rect 10048 44736 10100 44742
rect 10048 44678 10100 44684
rect 9109 44092 9417 44112
rect 9109 44090 9115 44092
rect 9171 44090 9195 44092
rect 9251 44090 9275 44092
rect 9331 44090 9355 44092
rect 9411 44090 9417 44092
rect 9171 44038 9173 44090
rect 9353 44038 9355 44090
rect 9109 44036 9115 44038
rect 9171 44036 9195 44038
rect 9251 44036 9275 44038
rect 9331 44036 9355 44038
rect 9411 44036 9417 44038
rect 9109 44016 9417 44036
rect 9876 43790 9904 44678
rect 10060 44441 10088 44678
rect 10046 44432 10102 44441
rect 10046 44367 10102 44376
rect 9864 43784 9916 43790
rect 9864 43726 9916 43732
rect 10046 43752 10102 43761
rect 10046 43687 10102 43696
rect 10060 43654 10088 43687
rect 9864 43648 9916 43654
rect 9864 43590 9916 43596
rect 10048 43648 10100 43654
rect 10048 43590 10100 43596
rect 9876 43314 9904 43590
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 10048 43104 10100 43110
rect 10048 43046 10100 43052
rect 9109 43004 9417 43024
rect 9109 43002 9115 43004
rect 9171 43002 9195 43004
rect 9251 43002 9275 43004
rect 9331 43002 9355 43004
rect 9411 43002 9417 43004
rect 9171 42950 9173 43002
rect 9353 42950 9355 43002
rect 9109 42948 9115 42950
rect 9171 42948 9195 42950
rect 9251 42948 9275 42950
rect 9331 42948 9355 42950
rect 9411 42948 9417 42950
rect 9109 42928 9417 42948
rect 10060 42945 10088 43046
rect 10046 42936 10102 42945
rect 10046 42871 10102 42880
rect 9864 42696 9916 42702
rect 9864 42638 9916 42644
rect 9109 41916 9417 41936
rect 9109 41914 9115 41916
rect 9171 41914 9195 41916
rect 9251 41914 9275 41916
rect 9331 41914 9355 41916
rect 9411 41914 9417 41916
rect 9171 41862 9173 41914
rect 9353 41862 9355 41914
rect 9109 41860 9115 41862
rect 9171 41860 9195 41862
rect 9251 41860 9275 41862
rect 9331 41860 9355 41862
rect 9411 41860 9417 41862
rect 9109 41840 9417 41860
rect 9876 41818 9904 42638
rect 10048 42560 10100 42566
rect 10048 42502 10100 42508
rect 10060 42265 10088 42502
rect 10046 42256 10102 42265
rect 10046 42191 10102 42200
rect 9864 41812 9916 41818
rect 9864 41754 9916 41760
rect 10048 41472 10100 41478
rect 10046 41440 10048 41449
rect 10100 41440 10102 41449
rect 10046 41375 10102 41384
rect 9864 41132 9916 41138
rect 9864 41074 9916 41080
rect 9109 40828 9417 40848
rect 9109 40826 9115 40828
rect 9171 40826 9195 40828
rect 9251 40826 9275 40828
rect 9331 40826 9355 40828
rect 9411 40826 9417 40828
rect 9171 40774 9173 40826
rect 9353 40774 9355 40826
rect 9109 40772 9115 40774
rect 9171 40772 9195 40774
rect 9251 40772 9275 40774
rect 9331 40772 9355 40774
rect 9411 40772 9417 40774
rect 9109 40752 9417 40772
rect 9109 39740 9417 39760
rect 9109 39738 9115 39740
rect 9171 39738 9195 39740
rect 9251 39738 9275 39740
rect 9331 39738 9355 39740
rect 9411 39738 9417 39740
rect 9171 39686 9173 39738
rect 9353 39686 9355 39738
rect 9109 39684 9115 39686
rect 9171 39684 9195 39686
rect 9251 39684 9275 39686
rect 9331 39684 9355 39686
rect 9411 39684 9417 39686
rect 9109 39664 9417 39684
rect 9876 39098 9904 41074
rect 10048 40928 10100 40934
rect 10048 40870 10100 40876
rect 10060 40633 10088 40870
rect 10046 40624 10102 40633
rect 10046 40559 10102 40568
rect 10046 39944 10102 39953
rect 10046 39879 10048 39888
rect 10100 39879 10102 39888
rect 10048 39850 10100 39856
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 10060 39137 10088 39238
rect 10046 39128 10102 39137
rect 9864 39092 9916 39098
rect 10046 39063 10102 39072
rect 9864 39034 9916 39040
rect 10048 38752 10100 38758
rect 10048 38694 10100 38700
rect 9109 38652 9417 38672
rect 9109 38650 9115 38652
rect 9171 38650 9195 38652
rect 9251 38650 9275 38652
rect 9331 38650 9355 38652
rect 9411 38650 9417 38652
rect 9171 38598 9173 38650
rect 9353 38598 9355 38650
rect 9109 38596 9115 38598
rect 9171 38596 9195 38598
rect 9251 38596 9275 38598
rect 9331 38596 9355 38598
rect 9411 38596 9417 38598
rect 9109 38576 9417 38596
rect 10060 38457 10088 38694
rect 10046 38448 10102 38457
rect 10046 38383 10102 38392
rect 9864 37868 9916 37874
rect 9864 37810 9916 37816
rect 9109 37564 9417 37584
rect 9109 37562 9115 37564
rect 9171 37562 9195 37564
rect 9251 37562 9275 37564
rect 9331 37562 9355 37564
rect 9411 37562 9417 37564
rect 9171 37510 9173 37562
rect 9353 37510 9355 37562
rect 9109 37508 9115 37510
rect 9171 37508 9195 37510
rect 9251 37508 9275 37510
rect 9331 37508 9355 37510
rect 9411 37508 9417 37510
rect 9109 37488 9417 37508
rect 9876 36922 9904 37810
rect 10048 37664 10100 37670
rect 10046 37632 10048 37641
rect 10100 37632 10102 37641
rect 10046 37567 10102 37576
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 9864 36916 9916 36922
rect 9864 36858 9916 36864
rect 10060 36825 10088 37062
rect 10046 36816 10102 36825
rect 10046 36751 10102 36760
rect 9109 36476 9417 36496
rect 9109 36474 9115 36476
rect 9171 36474 9195 36476
rect 9251 36474 9275 36476
rect 9331 36474 9355 36476
rect 9411 36474 9417 36476
rect 9171 36422 9173 36474
rect 9353 36422 9355 36474
rect 9109 36420 9115 36422
rect 9171 36420 9195 36422
rect 9251 36420 9275 36422
rect 9331 36420 9355 36422
rect 9411 36420 9417 36422
rect 9109 36400 9417 36420
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 10046 36136 10102 36145
rect 9772 35692 9824 35698
rect 9772 35634 9824 35640
rect 9109 35388 9417 35408
rect 9109 35386 9115 35388
rect 9171 35386 9195 35388
rect 9251 35386 9275 35388
rect 9331 35386 9355 35388
rect 9411 35386 9417 35388
rect 9171 35334 9173 35386
rect 9353 35334 9355 35386
rect 9109 35332 9115 35334
rect 9171 35332 9195 35334
rect 9251 35332 9275 35334
rect 9331 35332 9355 35334
rect 9411 35332 9417 35334
rect 9109 35312 9417 35332
rect 9784 35290 9812 35634
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9772 35080 9824 35086
rect 9772 35022 9824 35028
rect 9109 34300 9417 34320
rect 9109 34298 9115 34300
rect 9171 34298 9195 34300
rect 9251 34298 9275 34300
rect 9331 34298 9355 34300
rect 9411 34298 9417 34300
rect 9171 34246 9173 34298
rect 9353 34246 9355 34298
rect 9109 34244 9115 34246
rect 9171 34244 9195 34246
rect 9251 34244 9275 34246
rect 9331 34244 9355 34246
rect 9411 34244 9417 34246
rect 9109 34224 9417 34244
rect 9680 33992 9732 33998
rect 9680 33934 9732 33940
rect 9109 33212 9417 33232
rect 9109 33210 9115 33212
rect 9171 33210 9195 33212
rect 9251 33210 9275 33212
rect 9331 33210 9355 33212
rect 9411 33210 9417 33212
rect 9171 33158 9173 33210
rect 9353 33158 9355 33210
rect 9109 33156 9115 33158
rect 9171 33156 9195 33158
rect 9251 33156 9275 33158
rect 9331 33156 9355 33158
rect 9411 33156 9417 33158
rect 9109 33136 9417 33156
rect 9692 32570 9720 33934
rect 9784 33658 9812 35022
rect 9876 34202 9904 36110
rect 10046 36071 10102 36080
rect 10060 36038 10088 36071
rect 10048 36032 10100 36038
rect 10048 35974 10100 35980
rect 10048 35488 10100 35494
rect 10048 35430 10100 35436
rect 10060 35329 10088 35430
rect 10046 35320 10102 35329
rect 10046 35255 10102 35264
rect 10048 34944 10100 34950
rect 10048 34886 10100 34892
rect 10060 34649 10088 34886
rect 10046 34640 10102 34649
rect 10046 34575 10102 34584
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 10048 33856 10100 33862
rect 10046 33824 10048 33833
rect 10100 33824 10102 33833
rect 10046 33759 10102 33768
rect 9772 33652 9824 33658
rect 9772 33594 9824 33600
rect 9864 33516 9916 33522
rect 9864 33458 9916 33464
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9109 32124 9417 32144
rect 9109 32122 9115 32124
rect 9171 32122 9195 32124
rect 9251 32122 9275 32124
rect 9331 32122 9355 32124
rect 9411 32122 9417 32124
rect 9171 32070 9173 32122
rect 9353 32070 9355 32122
rect 9109 32068 9115 32070
rect 9171 32068 9195 32070
rect 9251 32068 9275 32070
rect 9331 32068 9355 32070
rect 9411 32068 9417 32070
rect 9109 32048 9417 32068
rect 9876 32026 9904 33458
rect 10048 33312 10100 33318
rect 10048 33254 10100 33260
rect 10060 33017 10088 33254
rect 10046 33008 10102 33017
rect 10046 32943 10102 32952
rect 10046 32328 10102 32337
rect 10046 32263 10048 32272
rect 10100 32263 10102 32272
rect 10048 32234 10100 32240
rect 9864 32020 9916 32026
rect 9864 31962 9916 31968
rect 10048 31680 10100 31686
rect 10048 31622 10100 31628
rect 10060 31521 10088 31622
rect 10046 31512 10102 31521
rect 10046 31447 10102 31456
rect 10048 31136 10100 31142
rect 10048 31078 10100 31084
rect 9109 31036 9417 31056
rect 9109 31034 9115 31036
rect 9171 31034 9195 31036
rect 9251 31034 9275 31036
rect 9331 31034 9355 31036
rect 9411 31034 9417 31036
rect 9171 30982 9173 31034
rect 9353 30982 9355 31034
rect 9109 30980 9115 30982
rect 9171 30980 9195 30982
rect 9251 30980 9275 30982
rect 9331 30980 9355 30982
rect 9411 30980 9417 30982
rect 9109 30960 9417 30980
rect 10060 30841 10088 31078
rect 10046 30832 10102 30841
rect 10046 30767 10102 30776
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 9109 29948 9417 29968
rect 9109 29946 9115 29948
rect 9171 29946 9195 29948
rect 9251 29946 9275 29948
rect 9331 29946 9355 29948
rect 9411 29946 9417 29948
rect 9171 29894 9173 29946
rect 9353 29894 9355 29946
rect 9109 29892 9115 29894
rect 9171 29892 9195 29894
rect 9251 29892 9275 29894
rect 9331 29892 9355 29894
rect 9411 29892 9417 29894
rect 9109 29872 9417 29892
rect 9109 28860 9417 28880
rect 9109 28858 9115 28860
rect 9171 28858 9195 28860
rect 9251 28858 9275 28860
rect 9331 28858 9355 28860
rect 9411 28858 9417 28860
rect 9171 28806 9173 28858
rect 9353 28806 9355 28858
rect 9109 28804 9115 28806
rect 9171 28804 9195 28806
rect 9251 28804 9275 28806
rect 9331 28804 9355 28806
rect 9411 28804 9417 28806
rect 9109 28784 9417 28804
rect 9109 27772 9417 27792
rect 9109 27770 9115 27772
rect 9171 27770 9195 27772
rect 9251 27770 9275 27772
rect 9331 27770 9355 27772
rect 9411 27770 9417 27772
rect 9171 27718 9173 27770
rect 9353 27718 9355 27770
rect 9109 27716 9115 27718
rect 9171 27716 9195 27718
rect 9251 27716 9275 27718
rect 9331 27716 9355 27718
rect 9411 27716 9417 27718
rect 9109 27696 9417 27716
rect 9876 27606 9904 30194
rect 10048 30048 10100 30054
rect 10046 30016 10048 30025
rect 10100 30016 10102 30025
rect 10046 29951 10102 29960
rect 10968 29232 11020 29238
rect 10966 29200 10968 29209
rect 11020 29200 11022 29209
rect 10966 29135 11022 29144
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28529 10180 28902
rect 10138 28520 10194 28529
rect 10138 28455 10194 28464
rect 10138 27704 10194 27713
rect 10138 27639 10140 27648
rect 10192 27639 10194 27648
rect 10140 27610 10192 27616
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 10138 27024 10194 27033
rect 10138 26959 10140 26968
rect 10192 26959 10194 26968
rect 10140 26930 10192 26936
rect 9109 26684 9417 26704
rect 9109 26682 9115 26684
rect 9171 26682 9195 26684
rect 9251 26682 9275 26684
rect 9331 26682 9355 26684
rect 9411 26682 9417 26684
rect 9171 26630 9173 26682
rect 9353 26630 9355 26682
rect 9109 26628 9115 26630
rect 9171 26628 9195 26630
rect 9251 26628 9275 26630
rect 9331 26628 9355 26630
rect 9411 26628 9417 26630
rect 9109 26608 9417 26628
rect 10138 26208 10194 26217
rect 10138 26143 10194 26152
rect 9109 25596 9417 25616
rect 9109 25594 9115 25596
rect 9171 25594 9195 25596
rect 9251 25594 9275 25596
rect 9331 25594 9355 25596
rect 9411 25594 9417 25596
rect 9171 25542 9173 25594
rect 9353 25542 9355 25594
rect 9109 25540 9115 25542
rect 9171 25540 9195 25542
rect 9251 25540 9275 25542
rect 9331 25540 9355 25542
rect 9411 25540 9417 25542
rect 9109 25520 9417 25540
rect 10152 25498 10180 26143
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10230 25392 10286 25401
rect 10230 25327 10286 25336
rect 10244 24886 10272 25327
rect 10232 24880 10284 24886
rect 10232 24822 10284 24828
rect 10138 24712 10194 24721
rect 10138 24647 10194 24656
rect 9109 24508 9417 24528
rect 9109 24506 9115 24508
rect 9171 24506 9195 24508
rect 9251 24506 9275 24508
rect 9331 24506 9355 24508
rect 9411 24506 9417 24508
rect 9171 24454 9173 24506
rect 9353 24454 9355 24506
rect 9109 24452 9115 24454
rect 9171 24452 9195 24454
rect 9251 24452 9275 24454
rect 9331 24452 9355 24454
rect 9411 24452 9417 24454
rect 9109 24432 9417 24452
rect 10152 24410 10180 24647
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10138 23896 10194 23905
rect 10138 23831 10194 23840
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9109 23420 9417 23440
rect 9109 23418 9115 23420
rect 9171 23418 9195 23420
rect 9251 23418 9275 23420
rect 9331 23418 9355 23420
rect 9411 23418 9417 23420
rect 9171 23366 9173 23418
rect 9353 23366 9355 23418
rect 9109 23364 9115 23366
rect 9171 23364 9195 23366
rect 9251 23364 9275 23366
rect 9331 23364 9355 23366
rect 9411 23364 9417 23366
rect 9109 23344 9417 23364
rect 9876 23322 9904 23666
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 10060 23225 10088 23462
rect 10152 23322 10180 23831
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10046 23216 10102 23225
rect 10046 23151 10102 23160
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 9109 22332 9417 22352
rect 9109 22330 9115 22332
rect 9171 22330 9195 22332
rect 9251 22330 9275 22332
rect 9331 22330 9355 22332
rect 9411 22330 9417 22332
rect 9171 22278 9173 22330
rect 9353 22278 9355 22330
rect 9109 22276 9115 22278
rect 9171 22276 9195 22278
rect 9251 22276 9275 22278
rect 9331 22276 9355 22278
rect 9411 22276 9417 22278
rect 9109 22256 9417 22276
rect 9109 21244 9417 21264
rect 9109 21242 9115 21244
rect 9171 21242 9195 21244
rect 9251 21242 9275 21244
rect 9331 21242 9355 21244
rect 9411 21242 9417 21244
rect 9171 21190 9173 21242
rect 9353 21190 9355 21242
rect 9109 21188 9115 21190
rect 9171 21188 9195 21190
rect 9251 21188 9275 21190
rect 9331 21188 9355 21190
rect 9411 21188 9417 21190
rect 9109 21168 9417 21188
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9109 20156 9417 20176
rect 9109 20154 9115 20156
rect 9171 20154 9195 20156
rect 9251 20154 9275 20156
rect 9331 20154 9355 20156
rect 9411 20154 9417 20156
rect 9171 20102 9173 20154
rect 9353 20102 9355 20154
rect 9109 20100 9115 20102
rect 9171 20100 9195 20102
rect 9251 20100 9275 20102
rect 9331 20100 9355 20102
rect 9411 20100 9417 20102
rect 9109 20080 9417 20100
rect 9109 19068 9417 19088
rect 9109 19066 9115 19068
rect 9171 19066 9195 19068
rect 9251 19066 9275 19068
rect 9331 19066 9355 19068
rect 9411 19066 9417 19068
rect 9171 19014 9173 19066
rect 9353 19014 9355 19066
rect 9109 19012 9115 19014
rect 9171 19012 9195 19014
rect 9251 19012 9275 19014
rect 9331 19012 9355 19014
rect 9411 19012 9417 19014
rect 9109 18992 9417 19012
rect 9784 18970 9812 20878
rect 9876 20602 9904 22578
rect 10048 22432 10100 22438
rect 10046 22400 10048 22409
rect 10100 22400 10102 22409
rect 10046 22335 10102 22344
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9109 17980 9417 18000
rect 9109 17978 9115 17980
rect 9171 17978 9195 17980
rect 9251 17978 9275 17980
rect 9331 17978 9355 17980
rect 9411 17978 9417 17980
rect 9171 17926 9173 17978
rect 9353 17926 9355 17978
rect 9109 17924 9115 17926
rect 9171 17924 9195 17926
rect 9251 17924 9275 17926
rect 9331 17924 9355 17926
rect 9411 17924 9417 17926
rect 9109 17904 9417 17924
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 9109 16892 9417 16912
rect 9109 16890 9115 16892
rect 9171 16890 9195 16892
rect 9251 16890 9275 16892
rect 9331 16890 9355 16892
rect 9411 16890 9417 16892
rect 9171 16838 9173 16890
rect 9353 16838 9355 16890
rect 9109 16836 9115 16838
rect 9171 16836 9195 16838
rect 9251 16836 9275 16838
rect 9331 16836 9355 16838
rect 9411 16836 9417 16838
rect 9109 16816 9417 16836
rect 9109 15804 9417 15824
rect 9109 15802 9115 15804
rect 9171 15802 9195 15804
rect 9251 15802 9275 15804
rect 9331 15802 9355 15804
rect 9411 15802 9417 15804
rect 9171 15750 9173 15802
rect 9353 15750 9355 15802
rect 9109 15748 9115 15750
rect 9171 15748 9195 15750
rect 9251 15748 9275 15750
rect 9331 15748 9355 15750
rect 9411 15748 9417 15750
rect 9109 15728 9417 15748
rect 9692 15570 9720 17614
rect 9784 16454 9812 18226
rect 9876 17882 9904 20402
rect 9968 19514 9996 21966
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21593 10088 21830
rect 10046 21584 10102 21593
rect 10046 21519 10102 21528
rect 10046 20904 10102 20913
rect 10046 20839 10102 20848
rect 10060 20806 10088 20839
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10060 20097 10088 20198
rect 10046 20088 10102 20097
rect 10046 20023 10102 20032
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10060 19417 10088 19654
rect 10046 19408 10102 19417
rect 10046 19343 10102 19352
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9876 15162 9904 16526
rect 9968 15706 9996 18702
rect 10048 18624 10100 18630
rect 10046 18592 10048 18601
rect 10100 18592 10102 18601
rect 10046 18527 10102 18536
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10060 17785 10088 18022
rect 10046 17776 10102 17785
rect 10046 17711 10102 17720
rect 10152 17270 10180 19314
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 10046 17096 10102 17105
rect 10046 17031 10048 17040
rect 10100 17031 10102 17040
rect 10048 17002 10100 17008
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16289 10088 16390
rect 10046 16280 10102 16289
rect 10046 16215 10102 16224
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10060 15609 10088 15846
rect 10046 15600 10102 15609
rect 10046 15535 10102 15544
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9864 15156 9916 15162
rect 9864 15098 9916 15104
rect 10048 14816 10100 14822
rect 10046 14784 10048 14793
rect 10100 14784 10102 14793
rect 9109 14716 9417 14736
rect 10046 14719 10102 14728
rect 9109 14714 9115 14716
rect 9171 14714 9195 14716
rect 9251 14714 9275 14716
rect 9331 14714 9355 14716
rect 9411 14714 9417 14716
rect 9171 14662 9173 14714
rect 9353 14662 9355 14714
rect 9109 14660 9115 14662
rect 9171 14660 9195 14662
rect 9251 14660 9275 14662
rect 9331 14660 9355 14662
rect 9411 14660 9417 14662
rect 9109 14640 9417 14660
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9109 13628 9417 13648
rect 9109 13626 9115 13628
rect 9171 13626 9195 13628
rect 9251 13626 9275 13628
rect 9331 13626 9355 13628
rect 9411 13626 9417 13628
rect 9171 13574 9173 13626
rect 9353 13574 9355 13626
rect 9109 13572 9115 13574
rect 9171 13572 9195 13574
rect 9251 13572 9275 13574
rect 9331 13572 9355 13574
rect 9411 13572 9417 13574
rect 9109 13552 9417 13572
rect 9109 12540 9417 12560
rect 9109 12538 9115 12540
rect 9171 12538 9195 12540
rect 9251 12538 9275 12540
rect 9331 12538 9355 12540
rect 9411 12538 9417 12540
rect 9171 12486 9173 12538
rect 9353 12486 9355 12538
rect 9109 12484 9115 12486
rect 9171 12484 9195 12486
rect 9251 12484 9275 12486
rect 9331 12484 9355 12486
rect 9411 12484 9417 12486
rect 9109 12464 9417 12484
rect 9784 12238 9812 13942
rect 9876 12850 9904 14010
rect 10060 13977 10088 14214
rect 10046 13968 10102 13977
rect 10046 13903 10102 13912
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 10046 13288 10102 13297
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9968 11898 9996 13262
rect 10046 13223 10102 13232
rect 10060 13190 10088 13223
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12481 10088 12582
rect 10046 12472 10102 12481
rect 10046 12407 10102 12416
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10060 11801 10088 12038
rect 10046 11792 10102 11801
rect 10046 11727 10102 11736
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9109 11452 9417 11472
rect 9109 11450 9115 11452
rect 9171 11450 9195 11452
rect 9251 11450 9275 11452
rect 9331 11450 9355 11452
rect 9411 11450 9417 11452
rect 9171 11398 9173 11450
rect 9353 11398 9355 11450
rect 9109 11396 9115 11398
rect 9171 11396 9195 11398
rect 9251 11396 9275 11398
rect 9331 11396 9355 11398
rect 9411 11396 9417 11398
rect 9109 11376 9417 11396
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 10048 11008 10100 11014
rect 10046 10976 10048 10985
rect 10100 10976 10102 10985
rect 10046 10911 10102 10920
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9109 10364 9417 10384
rect 9109 10362 9115 10364
rect 9171 10362 9195 10364
rect 9251 10362 9275 10364
rect 9331 10362 9355 10364
rect 9411 10362 9417 10364
rect 9171 10310 9173 10362
rect 9353 10310 9355 10362
rect 9109 10308 9115 10310
rect 9171 10308 9195 10310
rect 9251 10308 9275 10310
rect 9331 10308 9355 10310
rect 9411 10308 9417 10310
rect 9109 10288 9417 10308
rect 10060 10169 10088 10406
rect 10046 10160 10102 10169
rect 10046 10095 10102 10104
rect 10152 9654 10180 11698
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8404 8906 8432 9522
rect 10046 9480 10102 9489
rect 10046 9415 10048 9424
rect 10100 9415 10102 9424
rect 10048 9386 10100 9392
rect 9109 9276 9417 9296
rect 9109 9274 9115 9276
rect 9171 9274 9195 9276
rect 9251 9274 9275 9276
rect 9331 9274 9355 9276
rect 9411 9274 9417 9276
rect 9171 9222 9173 9274
rect 9353 9222 9355 9274
rect 9109 9220 9115 9222
rect 9171 9220 9195 9222
rect 9251 9220 9275 9222
rect 9331 9220 9355 9222
rect 9411 9220 9417 9222
rect 9109 9200 9417 9220
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9232 8498 9260 8774
rect 10060 8673 10088 8774
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9109 8188 9417 8208
rect 9109 8186 9115 8188
rect 9171 8186 9195 8188
rect 9251 8186 9275 8188
rect 9331 8186 9355 8188
rect 9411 8186 9417 8188
rect 9171 8134 9173 8186
rect 9353 8134 9355 8186
rect 9109 8132 9115 8134
rect 9171 8132 9195 8134
rect 9251 8132 9275 8134
rect 9331 8132 9355 8134
rect 9411 8132 9417 8134
rect 9109 8112 9417 8132
rect 10060 7993 10088 8230
rect 10046 7984 10102 7993
rect 10046 7919 10102 7928
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 7477 3292 7785 3312
rect 7477 3290 7483 3292
rect 7539 3290 7563 3292
rect 7619 3290 7643 3292
rect 7699 3290 7723 3292
rect 7779 3290 7785 3292
rect 7539 3238 7541 3290
rect 7721 3238 7723 3290
rect 7477 3236 7483 3238
rect 7539 3236 7563 3238
rect 7619 3236 7643 3238
rect 7699 3236 7723 3238
rect 7779 3236 7785 3238
rect 7477 3216 7785 3236
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5845 2748 6153 2768
rect 5845 2746 5851 2748
rect 5907 2746 5931 2748
rect 5987 2746 6011 2748
rect 6067 2746 6091 2748
rect 6147 2746 6153 2748
rect 5907 2694 5909 2746
rect 6089 2694 6091 2746
rect 5845 2692 5851 2694
rect 5907 2692 5931 2694
rect 5987 2692 6011 2694
rect 6067 2692 6091 2694
rect 6147 2692 6153 2694
rect 5845 2672 6153 2692
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 9048 2446 9076 7686
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9109 7100 9417 7120
rect 9109 7098 9115 7100
rect 9171 7098 9195 7100
rect 9251 7098 9275 7100
rect 9331 7098 9355 7100
rect 9411 7098 9417 7100
rect 9171 7046 9173 7098
rect 9353 7046 9355 7098
rect 9109 7044 9115 7046
rect 9171 7044 9195 7046
rect 9251 7044 9275 7046
rect 9331 7044 9355 7046
rect 9411 7044 9417 7046
rect 9109 7024 9417 7044
rect 9109 6012 9417 6032
rect 9109 6010 9115 6012
rect 9171 6010 9195 6012
rect 9251 6010 9275 6012
rect 9331 6010 9355 6012
rect 9411 6010 9417 6012
rect 9171 5958 9173 6010
rect 9353 5958 9355 6010
rect 9109 5956 9115 5958
rect 9171 5956 9195 5958
rect 9251 5956 9275 5958
rect 9331 5956 9355 5958
rect 9411 5956 9417 5958
rect 9109 5936 9417 5956
rect 9692 5846 9720 7346
rect 10048 7200 10100 7206
rect 10046 7168 10048 7177
rect 10100 7168 10102 7177
rect 10046 7103 10102 7112
rect 9772 6996 9824 7002
rect 9772 6938 9824 6944
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9109 4924 9417 4944
rect 9109 4922 9115 4924
rect 9171 4922 9195 4924
rect 9251 4922 9275 4924
rect 9331 4922 9355 4924
rect 9411 4922 9417 4924
rect 9171 4870 9173 4922
rect 9353 4870 9355 4922
rect 9109 4868 9115 4870
rect 9171 4868 9195 4870
rect 9251 4868 9275 4870
rect 9331 4868 9355 4870
rect 9411 4868 9417 4870
rect 9109 4848 9417 4868
rect 9692 4554 9720 5646
rect 9784 4622 9812 6938
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 6186 9904 6734
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6361 10088 6598
rect 10046 6352 10102 6361
rect 10046 6287 10102 6296
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 10046 5672 10102 5681
rect 10046 5607 10102 5616
rect 10060 5574 10088 5607
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4865 10088 4966
rect 10046 4856 10102 4865
rect 10046 4791 10102 4800
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9109 3836 9417 3856
rect 9109 3834 9115 3836
rect 9171 3834 9195 3836
rect 9251 3834 9275 3836
rect 9331 3834 9355 3836
rect 9411 3834 9417 3836
rect 9171 3782 9173 3834
rect 9353 3782 9355 3834
rect 9109 3780 9115 3782
rect 9171 3780 9195 3782
rect 9251 3780 9275 3782
rect 9331 3780 9355 3782
rect 9411 3780 9417 3782
rect 9109 3760 9417 3780
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9109 2748 9417 2768
rect 9109 2746 9115 2748
rect 9171 2746 9195 2748
rect 9251 2746 9275 2748
rect 9331 2746 9355 2748
rect 9411 2746 9417 2748
rect 9171 2694 9173 2746
rect 9353 2694 9355 2746
rect 9109 2692 9115 2694
rect 9171 2692 9195 2694
rect 9251 2692 9275 2694
rect 9331 2692 9355 2694
rect 9411 2692 9417 2694
rect 9109 2672 9417 2692
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 3988 1873 4016 2382
rect 4213 2204 4521 2224
rect 4213 2202 4219 2204
rect 4275 2202 4299 2204
rect 4355 2202 4379 2204
rect 4435 2202 4459 2204
rect 4515 2202 4521 2204
rect 4275 2150 4277 2202
rect 4457 2150 4459 2202
rect 4213 2148 4219 2150
rect 4275 2148 4299 2150
rect 4355 2148 4379 2150
rect 4435 2148 4459 2150
rect 4515 2148 4521 2150
rect 4213 2128 4521 2148
rect 3974 1864 4030 1873
rect 3974 1799 4030 1808
rect 3606 1048 3662 1057
rect 3606 983 3662 992
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 4632 542 4660 2382
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 7477 2204 7785 2224
rect 7477 2202 7483 2204
rect 7539 2202 7563 2204
rect 7619 2202 7643 2204
rect 7699 2202 7723 2204
rect 7779 2202 7785 2204
rect 7539 2150 7541 2202
rect 7721 2150 7723 2202
rect 7477 2148 7483 2150
rect 7539 2148 7563 2150
rect 7619 2148 7643 2150
rect 7699 2148 7723 2150
rect 7779 2148 7785 2150
rect 7477 2128 7785 2148
rect 2780 536 2832 542
rect 2780 478 2832 484
rect 4620 536 4672 542
rect 4620 478 4672 484
rect 2792 241 2820 478
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 5998 0 6054 800
rect 9324 377 9352 2246
rect 9508 1873 9536 2790
rect 9784 2446 9812 4218
rect 10060 4185 10088 4422
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9876 3058 9904 3946
rect 10048 3392 10100 3398
rect 10046 3360 10048 3369
rect 10100 3360 10102 3369
rect 10046 3295 10102 3304
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2553 10088 2790
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 9494 1864 9550 1873
rect 9494 1799 9550 1808
rect 10060 1057 10088 2246
rect 10046 1048 10102 1057
rect 10046 983 10102 992
rect 9310 368 9366 377
rect 9310 303 9366 312
<< via2 >>
rect 2962 79600 3018 79656
rect 2588 77818 2644 77820
rect 2668 77818 2724 77820
rect 2748 77818 2804 77820
rect 2828 77818 2884 77820
rect 2588 77766 2634 77818
rect 2634 77766 2644 77818
rect 2668 77766 2698 77818
rect 2698 77766 2710 77818
rect 2710 77766 2724 77818
rect 2748 77766 2762 77818
rect 2762 77766 2774 77818
rect 2774 77766 2804 77818
rect 2828 77766 2838 77818
rect 2838 77766 2884 77818
rect 2588 77764 2644 77766
rect 2668 77764 2724 77766
rect 2748 77764 2804 77766
rect 2828 77764 2884 77766
rect 846 58792 902 58848
rect 3882 79192 3938 79248
rect 3054 78784 3110 78840
rect 3330 78376 3386 78432
rect 2502 77016 2558 77072
rect 1122 57468 1124 57488
rect 1124 57468 1176 57488
rect 1176 57468 1178 57488
rect 1122 57432 1178 57468
rect 1398 75384 1454 75440
rect 1306 74024 1362 74080
rect 2778 76880 2834 76936
rect 2042 76200 2098 76256
rect 1398 73616 1454 73672
rect 1398 72392 1454 72448
rect 1306 71848 1362 71904
rect 1306 71440 1362 71496
rect 1398 71032 1454 71088
rect 1306 70216 1362 70272
rect 1582 69672 1638 69728
rect 1766 72120 1822 72176
rect 1766 69436 1768 69456
rect 1768 69436 1820 69456
rect 1820 69436 1822 69456
rect 1766 69400 1822 69436
rect 1490 68992 1546 69048
rect 1306 67632 1362 67688
rect 1398 67224 1454 67280
rect 1398 65864 1454 65920
rect 1490 65456 1546 65512
rect 1490 64232 1546 64288
rect 1398 62464 1454 62520
rect 1490 61648 1546 61704
rect 2588 76730 2644 76732
rect 2668 76730 2724 76732
rect 2748 76730 2804 76732
rect 2828 76730 2884 76732
rect 2588 76678 2634 76730
rect 2634 76678 2644 76730
rect 2668 76678 2698 76730
rect 2698 76678 2710 76730
rect 2710 76678 2724 76730
rect 2748 76678 2762 76730
rect 2762 76678 2774 76730
rect 2774 76678 2804 76730
rect 2828 76678 2838 76730
rect 2838 76678 2884 76730
rect 2588 76676 2644 76678
rect 2668 76676 2724 76678
rect 2748 76676 2804 76678
rect 2828 76676 2884 76678
rect 2962 75792 3018 75848
rect 2588 75642 2644 75644
rect 2668 75642 2724 75644
rect 2748 75642 2804 75644
rect 2828 75642 2884 75644
rect 2588 75590 2634 75642
rect 2634 75590 2644 75642
rect 2668 75590 2698 75642
rect 2698 75590 2710 75642
rect 2710 75590 2724 75642
rect 2748 75590 2762 75642
rect 2762 75590 2774 75642
rect 2774 75590 2804 75642
rect 2828 75590 2838 75642
rect 2838 75590 2884 75642
rect 2588 75588 2644 75590
rect 2668 75588 2724 75590
rect 2748 75588 2804 75590
rect 2828 75588 2884 75590
rect 2588 74554 2644 74556
rect 2668 74554 2724 74556
rect 2748 74554 2804 74556
rect 2828 74554 2884 74556
rect 2588 74502 2634 74554
rect 2634 74502 2644 74554
rect 2668 74502 2698 74554
rect 2698 74502 2710 74554
rect 2710 74502 2724 74554
rect 2748 74502 2762 74554
rect 2762 74502 2774 74554
rect 2774 74502 2804 74554
rect 2828 74502 2838 74554
rect 2838 74502 2884 74554
rect 2588 74500 2644 74502
rect 2668 74500 2724 74502
rect 2748 74500 2804 74502
rect 2828 74500 2884 74502
rect 2226 72800 2282 72856
rect 2134 72120 2190 72176
rect 1490 59880 1546 59936
rect 1398 59508 1400 59528
rect 1400 59508 1452 59528
rect 1452 59508 1454 59528
rect 1398 59472 1454 59508
rect 1306 59064 1362 59120
rect 1306 57840 1362 57896
rect 1490 58112 1546 58168
rect 1398 57296 1454 57352
rect 1398 56888 1454 56944
rect 1490 56480 1546 56536
rect 1490 54712 1546 54768
rect 1490 53896 1546 53952
rect 1398 52128 1454 52184
rect 1490 51720 1546 51776
rect 1306 51032 1362 51088
rect 1306 50496 1362 50552
rect 2042 61920 2098 61976
rect 1858 57840 1914 57896
rect 2588 73466 2644 73468
rect 2668 73466 2724 73468
rect 2748 73466 2804 73468
rect 2828 73466 2884 73468
rect 2588 73414 2634 73466
rect 2634 73414 2644 73466
rect 2668 73414 2698 73466
rect 2698 73414 2710 73466
rect 2710 73414 2724 73466
rect 2748 73414 2762 73466
rect 2762 73414 2774 73466
rect 2774 73414 2804 73466
rect 2828 73414 2838 73466
rect 2838 73414 2884 73466
rect 2588 73412 2644 73414
rect 2668 73412 2724 73414
rect 2748 73412 2804 73414
rect 2828 73412 2884 73414
rect 2962 73208 3018 73264
rect 2588 72378 2644 72380
rect 2668 72378 2724 72380
rect 2748 72378 2804 72380
rect 2828 72378 2884 72380
rect 2588 72326 2634 72378
rect 2634 72326 2644 72378
rect 2668 72326 2698 72378
rect 2698 72326 2710 72378
rect 2710 72326 2724 72378
rect 2748 72326 2762 72378
rect 2762 72326 2774 72378
rect 2774 72326 2804 72378
rect 2828 72326 2838 72378
rect 2838 72326 2884 72378
rect 2588 72324 2644 72326
rect 2668 72324 2724 72326
rect 2748 72324 2804 72326
rect 2828 72324 2884 72326
rect 2588 71290 2644 71292
rect 2668 71290 2724 71292
rect 2748 71290 2804 71292
rect 2828 71290 2884 71292
rect 2588 71238 2634 71290
rect 2634 71238 2644 71290
rect 2668 71238 2698 71290
rect 2698 71238 2710 71290
rect 2710 71238 2724 71290
rect 2748 71238 2762 71290
rect 2762 71238 2774 71290
rect 2774 71238 2804 71290
rect 2828 71238 2838 71290
rect 2838 71238 2884 71290
rect 2588 71236 2644 71238
rect 2668 71236 2724 71238
rect 2748 71236 2804 71238
rect 2828 71236 2884 71238
rect 2410 69672 2466 69728
rect 2318 66272 2374 66328
rect 2318 64776 2374 64832
rect 2226 62056 2282 62112
rect 2226 61920 2282 61976
rect 1490 49952 1546 50008
rect 2778 70624 2834 70680
rect 2588 70202 2644 70204
rect 2668 70202 2724 70204
rect 2748 70202 2804 70204
rect 2828 70202 2884 70204
rect 2588 70150 2634 70202
rect 2634 70150 2644 70202
rect 2668 70150 2698 70202
rect 2698 70150 2710 70202
rect 2710 70150 2724 70202
rect 2748 70150 2762 70202
rect 2762 70150 2774 70202
rect 2774 70150 2804 70202
rect 2828 70150 2838 70202
rect 2838 70150 2884 70202
rect 2588 70148 2644 70150
rect 2668 70148 2724 70150
rect 2748 70148 2804 70150
rect 2828 70148 2884 70150
rect 10138 78648 10194 78704
rect 4066 77968 4122 78024
rect 3974 77560 4030 77616
rect 5851 77818 5907 77820
rect 5931 77818 5987 77820
rect 6011 77818 6067 77820
rect 6091 77818 6147 77820
rect 5851 77766 5897 77818
rect 5897 77766 5907 77818
rect 5931 77766 5961 77818
rect 5961 77766 5973 77818
rect 5973 77766 5987 77818
rect 6011 77766 6025 77818
rect 6025 77766 6037 77818
rect 6037 77766 6067 77818
rect 6091 77766 6101 77818
rect 6101 77766 6147 77818
rect 5851 77764 5907 77766
rect 5931 77764 5987 77766
rect 6011 77764 6067 77766
rect 6091 77764 6147 77766
rect 9115 77818 9171 77820
rect 9195 77818 9251 77820
rect 9275 77818 9331 77820
rect 9355 77818 9411 77820
rect 9115 77766 9161 77818
rect 9161 77766 9171 77818
rect 9195 77766 9225 77818
rect 9225 77766 9237 77818
rect 9237 77766 9251 77818
rect 9275 77766 9289 77818
rect 9289 77766 9301 77818
rect 9301 77766 9331 77818
rect 9355 77766 9365 77818
rect 9365 77766 9411 77818
rect 9115 77764 9171 77766
rect 9195 77764 9251 77766
rect 9275 77764 9331 77766
rect 9355 77764 9411 77766
rect 4219 77274 4275 77276
rect 4299 77274 4355 77276
rect 4379 77274 4435 77276
rect 4459 77274 4515 77276
rect 4219 77222 4265 77274
rect 4265 77222 4275 77274
rect 4299 77222 4329 77274
rect 4329 77222 4341 77274
rect 4341 77222 4355 77274
rect 4379 77222 4393 77274
rect 4393 77222 4405 77274
rect 4405 77222 4435 77274
rect 4459 77222 4469 77274
rect 4469 77222 4515 77274
rect 4219 77220 4275 77222
rect 4299 77220 4355 77222
rect 4379 77220 4435 77222
rect 4459 77220 4515 77222
rect 3606 74296 3662 74352
rect 4219 76186 4275 76188
rect 4299 76186 4355 76188
rect 4379 76186 4435 76188
rect 4459 76186 4515 76188
rect 4219 76134 4265 76186
rect 4265 76134 4275 76186
rect 4299 76134 4329 76186
rect 4329 76134 4341 76186
rect 4341 76134 4355 76186
rect 4379 76134 4393 76186
rect 4393 76134 4405 76186
rect 4405 76134 4435 76186
rect 4459 76134 4469 76186
rect 4469 76134 4515 76186
rect 4219 76132 4275 76134
rect 4299 76132 4355 76134
rect 4379 76132 4435 76134
rect 4459 76132 4515 76134
rect 4219 75098 4275 75100
rect 4299 75098 4355 75100
rect 4379 75098 4435 75100
rect 4459 75098 4515 75100
rect 4219 75046 4265 75098
rect 4265 75046 4275 75098
rect 4299 75046 4329 75098
rect 4329 75046 4341 75098
rect 4341 75046 4355 75098
rect 4379 75046 4393 75098
rect 4393 75046 4405 75098
rect 4405 75046 4435 75098
rect 4459 75046 4469 75098
rect 4469 75046 4515 75098
rect 4219 75044 4275 75046
rect 4299 75044 4355 75046
rect 4379 75044 4435 75046
rect 4459 75044 4515 75046
rect 3974 74976 4030 75032
rect 10966 77988 11022 78024
rect 10966 77968 10968 77988
rect 10968 77968 11020 77988
rect 11020 77968 11022 77988
rect 7483 77274 7539 77276
rect 7563 77274 7619 77276
rect 7643 77274 7699 77276
rect 7723 77274 7779 77276
rect 7483 77222 7529 77274
rect 7529 77222 7539 77274
rect 7563 77222 7593 77274
rect 7593 77222 7605 77274
rect 7605 77222 7619 77274
rect 7643 77222 7657 77274
rect 7657 77222 7669 77274
rect 7669 77222 7699 77274
rect 7723 77222 7733 77274
rect 7733 77222 7779 77274
rect 7483 77220 7539 77222
rect 7563 77220 7619 77222
rect 7643 77220 7699 77222
rect 7723 77220 7779 77222
rect 9402 77152 9458 77208
rect 5851 76730 5907 76732
rect 5931 76730 5987 76732
rect 6011 76730 6067 76732
rect 6091 76730 6147 76732
rect 5851 76678 5897 76730
rect 5897 76678 5907 76730
rect 5931 76678 5961 76730
rect 5961 76678 5973 76730
rect 5973 76678 5987 76730
rect 6011 76678 6025 76730
rect 6025 76678 6037 76730
rect 6037 76678 6067 76730
rect 6091 76678 6101 76730
rect 6101 76678 6147 76730
rect 5851 76676 5907 76678
rect 5931 76676 5987 76678
rect 6011 76676 6067 76678
rect 6091 76676 6147 76678
rect 9115 76730 9171 76732
rect 9195 76730 9251 76732
rect 9275 76730 9331 76732
rect 9355 76730 9411 76732
rect 9115 76678 9161 76730
rect 9161 76678 9171 76730
rect 9195 76678 9225 76730
rect 9225 76678 9237 76730
rect 9237 76678 9251 76730
rect 9275 76678 9289 76730
rect 9289 76678 9301 76730
rect 9301 76678 9331 76730
rect 9355 76678 9365 76730
rect 9365 76678 9411 76730
rect 9115 76676 9171 76678
rect 9195 76676 9251 76678
rect 9275 76676 9331 76678
rect 9355 76676 9411 76678
rect 7483 76186 7539 76188
rect 7563 76186 7619 76188
rect 7643 76186 7699 76188
rect 7723 76186 7779 76188
rect 7483 76134 7529 76186
rect 7529 76134 7539 76186
rect 7563 76134 7593 76186
rect 7593 76134 7605 76186
rect 7605 76134 7619 76186
rect 7643 76134 7657 76186
rect 7657 76134 7669 76186
rect 7669 76134 7699 76186
rect 7723 76134 7733 76186
rect 7733 76134 7779 76186
rect 7483 76132 7539 76134
rect 7563 76132 7619 76134
rect 7643 76132 7699 76134
rect 7723 76132 7779 76134
rect 5851 75642 5907 75644
rect 5931 75642 5987 75644
rect 6011 75642 6067 75644
rect 6091 75642 6147 75644
rect 5851 75590 5897 75642
rect 5897 75590 5907 75642
rect 5931 75590 5961 75642
rect 5961 75590 5973 75642
rect 5973 75590 5987 75642
rect 6011 75590 6025 75642
rect 6025 75590 6037 75642
rect 6037 75590 6067 75642
rect 6091 75590 6101 75642
rect 6101 75590 6147 75642
rect 5851 75588 5907 75590
rect 5931 75588 5987 75590
rect 6011 75588 6067 75590
rect 6091 75588 6147 75590
rect 3514 69808 3570 69864
rect 2588 69114 2644 69116
rect 2668 69114 2724 69116
rect 2748 69114 2804 69116
rect 2828 69114 2884 69116
rect 2588 69062 2634 69114
rect 2634 69062 2644 69114
rect 2668 69062 2698 69114
rect 2698 69062 2710 69114
rect 2710 69062 2724 69114
rect 2748 69062 2762 69114
rect 2762 69062 2774 69114
rect 2774 69062 2804 69114
rect 2828 69062 2838 69114
rect 2838 69062 2884 69114
rect 2588 69060 2644 69062
rect 2668 69060 2724 69062
rect 2748 69060 2804 69062
rect 2828 69060 2884 69062
rect 2588 68026 2644 68028
rect 2668 68026 2724 68028
rect 2748 68026 2804 68028
rect 2828 68026 2884 68028
rect 2588 67974 2634 68026
rect 2634 67974 2644 68026
rect 2668 67974 2698 68026
rect 2698 67974 2710 68026
rect 2710 67974 2724 68026
rect 2748 67974 2762 68026
rect 2762 67974 2774 68026
rect 2774 67974 2804 68026
rect 2828 67974 2838 68026
rect 2838 67974 2884 68026
rect 2588 67972 2644 67974
rect 2668 67972 2724 67974
rect 2748 67972 2804 67974
rect 2828 67972 2884 67974
rect 2588 66938 2644 66940
rect 2668 66938 2724 66940
rect 2748 66938 2804 66940
rect 2828 66938 2884 66940
rect 2588 66886 2634 66938
rect 2634 66886 2644 66938
rect 2668 66886 2698 66938
rect 2698 66886 2710 66938
rect 2710 66886 2724 66938
rect 2748 66886 2762 66938
rect 2762 66886 2774 66938
rect 2774 66886 2804 66938
rect 2828 66886 2838 66938
rect 2838 66886 2884 66938
rect 2588 66884 2644 66886
rect 2668 66884 2724 66886
rect 2748 66884 2804 66886
rect 2828 66884 2884 66886
rect 2962 66680 3018 66736
rect 2588 65850 2644 65852
rect 2668 65850 2724 65852
rect 2748 65850 2804 65852
rect 2828 65850 2884 65852
rect 2588 65798 2634 65850
rect 2634 65798 2644 65850
rect 2668 65798 2698 65850
rect 2698 65798 2710 65850
rect 2710 65798 2724 65850
rect 2748 65798 2762 65850
rect 2762 65798 2774 65850
rect 2774 65798 2804 65850
rect 2828 65798 2838 65850
rect 2838 65798 2884 65850
rect 2588 65796 2644 65798
rect 2668 65796 2724 65798
rect 2748 65796 2804 65798
rect 2828 65796 2884 65798
rect 2588 64762 2644 64764
rect 2668 64762 2724 64764
rect 2748 64762 2804 64764
rect 2828 64762 2884 64764
rect 2588 64710 2634 64762
rect 2634 64710 2644 64762
rect 2668 64710 2698 64762
rect 2698 64710 2710 64762
rect 2710 64710 2724 64762
rect 2748 64710 2762 64762
rect 2762 64710 2774 64762
rect 2774 64710 2804 64762
rect 2828 64710 2838 64762
rect 2838 64710 2884 64762
rect 2588 64708 2644 64710
rect 2668 64708 2724 64710
rect 2748 64708 2804 64710
rect 2828 64708 2884 64710
rect 2588 63674 2644 63676
rect 2668 63674 2724 63676
rect 2748 63674 2804 63676
rect 2828 63674 2884 63676
rect 2588 63622 2634 63674
rect 2634 63622 2644 63674
rect 2668 63622 2698 63674
rect 2698 63622 2710 63674
rect 2710 63622 2724 63674
rect 2748 63622 2762 63674
rect 2762 63622 2774 63674
rect 2774 63622 2804 63674
rect 2828 63622 2838 63674
rect 2838 63622 2884 63674
rect 2588 63620 2644 63622
rect 2668 63620 2724 63622
rect 2748 63620 2804 63622
rect 2828 63620 2884 63622
rect 2870 63436 2926 63472
rect 2870 63416 2872 63436
rect 2872 63416 2924 63436
rect 2924 63416 2926 63436
rect 2870 63144 2926 63200
rect 2588 62586 2644 62588
rect 2668 62586 2724 62588
rect 2748 62586 2804 62588
rect 2828 62586 2884 62588
rect 2588 62534 2634 62586
rect 2634 62534 2644 62586
rect 2668 62534 2698 62586
rect 2698 62534 2710 62586
rect 2710 62534 2724 62586
rect 2748 62534 2762 62586
rect 2762 62534 2774 62586
rect 2774 62534 2804 62586
rect 2828 62534 2838 62586
rect 2838 62534 2884 62586
rect 2588 62532 2644 62534
rect 2668 62532 2724 62534
rect 2748 62532 2804 62534
rect 2828 62532 2884 62534
rect 3054 65048 3110 65104
rect 3146 63280 3202 63336
rect 2588 61498 2644 61500
rect 2668 61498 2724 61500
rect 2748 61498 2804 61500
rect 2828 61498 2884 61500
rect 2588 61446 2634 61498
rect 2634 61446 2644 61498
rect 2668 61446 2698 61498
rect 2698 61446 2710 61498
rect 2710 61446 2724 61498
rect 2748 61446 2762 61498
rect 2762 61446 2774 61498
rect 2774 61446 2804 61498
rect 2828 61446 2838 61498
rect 2838 61446 2884 61498
rect 2588 61444 2644 61446
rect 2668 61444 2724 61446
rect 2748 61444 2804 61446
rect 2828 61444 2884 61446
rect 2962 60696 3018 60752
rect 2778 60560 2834 60616
rect 2588 60410 2644 60412
rect 2668 60410 2724 60412
rect 2748 60410 2804 60412
rect 2828 60410 2884 60412
rect 2588 60358 2634 60410
rect 2634 60358 2644 60410
rect 2668 60358 2698 60410
rect 2698 60358 2710 60410
rect 2710 60358 2724 60410
rect 2748 60358 2762 60410
rect 2762 60358 2774 60410
rect 2774 60358 2804 60410
rect 2828 60358 2838 60410
rect 2838 60358 2884 60410
rect 2588 60356 2644 60358
rect 2668 60356 2724 60358
rect 2748 60356 2804 60358
rect 2828 60356 2884 60358
rect 2588 59322 2644 59324
rect 2668 59322 2724 59324
rect 2748 59322 2804 59324
rect 2828 59322 2884 59324
rect 2588 59270 2634 59322
rect 2634 59270 2644 59322
rect 2668 59270 2698 59322
rect 2698 59270 2710 59322
rect 2710 59270 2724 59322
rect 2748 59270 2762 59322
rect 2762 59270 2774 59322
rect 2774 59270 2804 59322
rect 2828 59270 2838 59322
rect 2838 59270 2884 59322
rect 2588 59268 2644 59270
rect 2668 59268 2724 59270
rect 2748 59268 2804 59270
rect 2828 59268 2884 59270
rect 2588 58234 2644 58236
rect 2668 58234 2724 58236
rect 2748 58234 2804 58236
rect 2828 58234 2884 58236
rect 2588 58182 2634 58234
rect 2634 58182 2644 58234
rect 2668 58182 2698 58234
rect 2698 58182 2710 58234
rect 2710 58182 2724 58234
rect 2748 58182 2762 58234
rect 2762 58182 2774 58234
rect 2774 58182 2804 58234
rect 2828 58182 2838 58234
rect 2838 58182 2884 58234
rect 2588 58180 2644 58182
rect 2668 58180 2724 58182
rect 2748 58180 2804 58182
rect 2828 58180 2884 58182
rect 2778 57740 2780 57760
rect 2780 57740 2832 57760
rect 2832 57740 2834 57760
rect 2778 57704 2834 57740
rect 2870 57296 2926 57352
rect 2588 57146 2644 57148
rect 2668 57146 2724 57148
rect 2748 57146 2804 57148
rect 2828 57146 2884 57148
rect 2588 57094 2634 57146
rect 2634 57094 2644 57146
rect 2668 57094 2698 57146
rect 2698 57094 2710 57146
rect 2710 57094 2724 57146
rect 2748 57094 2762 57146
rect 2762 57094 2774 57146
rect 2774 57094 2804 57146
rect 2828 57094 2838 57146
rect 2838 57094 2884 57146
rect 2588 57092 2644 57094
rect 2668 57092 2724 57094
rect 2748 57092 2804 57094
rect 2828 57092 2884 57094
rect 2226 54576 2282 54632
rect 2226 54304 2282 54360
rect 3422 68176 3478 68232
rect 3330 60696 3386 60752
rect 3238 57432 3294 57488
rect 3146 56208 3202 56264
rect 2588 56058 2644 56060
rect 2668 56058 2724 56060
rect 2748 56058 2804 56060
rect 2828 56058 2884 56060
rect 2588 56006 2634 56058
rect 2634 56006 2644 56058
rect 2668 56006 2698 56058
rect 2698 56006 2710 56058
rect 2710 56006 2724 56058
rect 2748 56006 2762 56058
rect 2762 56006 2774 56058
rect 2774 56006 2804 56058
rect 2828 56006 2838 56058
rect 2838 56006 2884 56058
rect 2588 56004 2644 56006
rect 2668 56004 2724 56006
rect 2748 56004 2804 56006
rect 2828 56004 2884 56006
rect 2778 55140 2834 55176
rect 2778 55120 2780 55140
rect 2780 55120 2832 55140
rect 2832 55120 2834 55140
rect 2588 54970 2644 54972
rect 2668 54970 2724 54972
rect 2748 54970 2804 54972
rect 2828 54970 2884 54972
rect 2588 54918 2634 54970
rect 2634 54918 2644 54970
rect 2668 54918 2698 54970
rect 2698 54918 2710 54970
rect 2710 54918 2724 54970
rect 2748 54918 2762 54970
rect 2762 54918 2774 54970
rect 2774 54918 2804 54970
rect 2828 54918 2838 54970
rect 2838 54918 2884 54970
rect 2588 54916 2644 54918
rect 2668 54916 2724 54918
rect 2748 54916 2804 54918
rect 2828 54916 2884 54918
rect 3146 55800 3202 55856
rect 3146 55392 3202 55448
rect 2588 53882 2644 53884
rect 2668 53882 2724 53884
rect 2748 53882 2804 53884
rect 2828 53882 2884 53884
rect 2588 53830 2634 53882
rect 2634 53830 2644 53882
rect 2668 53830 2698 53882
rect 2698 53830 2710 53882
rect 2710 53830 2724 53882
rect 2748 53830 2762 53882
rect 2762 53830 2774 53882
rect 2774 53830 2804 53882
rect 2828 53830 2838 53882
rect 2838 53830 2884 53882
rect 2588 53828 2644 53830
rect 2668 53828 2724 53830
rect 2748 53828 2804 53830
rect 2828 53828 2884 53830
rect 2778 53488 2834 53544
rect 2226 52536 2282 52592
rect 2226 51312 2282 51368
rect 2134 51176 2190 51232
rect 2226 50924 2282 50960
rect 2226 50904 2228 50924
rect 2228 50904 2280 50924
rect 2280 50904 2282 50924
rect 2134 50768 2190 50824
rect 2042 50632 2098 50688
rect 1490 48320 1546 48376
rect 1490 47776 1546 47832
rect 1490 46960 1546 47016
rect 1490 46552 1546 46608
rect 1490 46144 1546 46200
rect 1490 45228 1492 45248
rect 1492 45228 1544 45248
rect 1544 45228 1546 45248
rect 1490 45192 1546 45228
rect 1582 44376 1638 44432
rect 1490 42200 1546 42256
rect 1398 41792 1454 41848
rect 1490 41384 1546 41440
rect 1950 49000 2006 49056
rect 1858 42200 1914 42256
rect 2226 49136 2282 49192
rect 2226 48592 2282 48648
rect 2226 47404 2228 47424
rect 2228 47404 2280 47424
rect 2280 47404 2282 47424
rect 2226 47368 2282 47404
rect 2588 52794 2644 52796
rect 2668 52794 2724 52796
rect 2748 52794 2804 52796
rect 2828 52794 2884 52796
rect 2588 52742 2634 52794
rect 2634 52742 2644 52794
rect 2668 52742 2698 52794
rect 2698 52742 2710 52794
rect 2710 52742 2724 52794
rect 2748 52742 2762 52794
rect 2762 52742 2774 52794
rect 2774 52742 2804 52794
rect 2828 52742 2838 52794
rect 2838 52742 2884 52794
rect 2588 52740 2644 52742
rect 2668 52740 2724 52742
rect 2748 52740 2804 52742
rect 2828 52740 2884 52742
rect 3054 52964 3110 53000
rect 3054 52944 3056 52964
rect 3056 52944 3108 52964
rect 3108 52944 3110 52964
rect 2588 51706 2644 51708
rect 2668 51706 2724 51708
rect 2748 51706 2804 51708
rect 2828 51706 2884 51708
rect 2588 51654 2634 51706
rect 2634 51654 2644 51706
rect 2668 51654 2698 51706
rect 2698 51654 2710 51706
rect 2710 51654 2724 51706
rect 2748 51654 2762 51706
rect 2762 51654 2774 51706
rect 2774 51654 2804 51706
rect 2828 51654 2838 51706
rect 2838 51654 2884 51706
rect 2588 51652 2644 51654
rect 2668 51652 2724 51654
rect 2748 51652 2804 51654
rect 2828 51652 2884 51654
rect 2502 51040 2558 51096
rect 2502 50768 2558 50824
rect 2778 50924 2834 50960
rect 2778 50904 2780 50924
rect 2780 50904 2832 50924
rect 2832 50904 2834 50924
rect 2410 49680 2466 49736
rect 2410 49580 2412 49600
rect 2412 49580 2464 49600
rect 2464 49580 2466 49600
rect 2410 49544 2466 49580
rect 2134 46008 2190 46064
rect 2042 45056 2098 45112
rect 2318 46416 2374 46472
rect 2410 45600 2466 45656
rect 2410 44784 2466 44840
rect 2410 43968 2466 44024
rect 2318 43424 2374 43480
rect 2226 43152 2282 43208
rect 2226 42608 2282 42664
rect 1858 41792 1914 41848
rect 1766 41248 1822 41304
rect 1398 40568 1454 40624
rect 1490 39208 1546 39264
rect 1398 37984 1454 38040
rect 1674 41112 1730 41168
rect 1490 37032 1546 37088
rect 1490 36080 1546 36136
rect 1398 35808 1454 35864
rect 1398 35672 1454 35728
rect 1490 35400 1546 35456
rect 1490 34992 1546 35048
rect 1490 33224 1546 33280
rect 1398 32408 1454 32464
rect 1214 31864 1270 31920
rect 1214 24248 1270 24304
rect 1214 22072 1270 22128
rect 1214 15544 1270 15600
rect 1122 14728 1178 14784
rect 1490 30640 1546 30696
rect 1674 32000 1730 32056
rect 1766 31728 1822 31784
rect 1398 28056 1454 28112
rect 2042 42064 2098 42120
rect 2134 41248 2190 41304
rect 2318 41248 2374 41304
rect 2318 40996 2374 41032
rect 2318 40976 2320 40996
rect 2320 40976 2372 40996
rect 2372 40976 2374 40996
rect 2318 39616 2374 39672
rect 2870 50768 2926 50824
rect 2588 50618 2644 50620
rect 2668 50618 2724 50620
rect 2748 50618 2804 50620
rect 2828 50618 2884 50620
rect 2588 50566 2634 50618
rect 2634 50566 2644 50618
rect 2668 50566 2698 50618
rect 2698 50566 2710 50618
rect 2710 50566 2724 50618
rect 2748 50566 2762 50618
rect 2762 50566 2774 50618
rect 2774 50566 2804 50618
rect 2828 50566 2838 50618
rect 2838 50566 2884 50618
rect 2588 50564 2644 50566
rect 2668 50564 2724 50566
rect 2748 50564 2804 50566
rect 2828 50564 2884 50566
rect 2588 49530 2644 49532
rect 2668 49530 2724 49532
rect 2748 49530 2804 49532
rect 2828 49530 2884 49532
rect 2588 49478 2634 49530
rect 2634 49478 2644 49530
rect 2668 49478 2698 49530
rect 2698 49478 2710 49530
rect 2710 49478 2724 49530
rect 2748 49478 2762 49530
rect 2762 49478 2774 49530
rect 2774 49478 2804 49530
rect 2828 49478 2838 49530
rect 2838 49478 2884 49530
rect 2588 49476 2644 49478
rect 2668 49476 2724 49478
rect 2748 49476 2804 49478
rect 2828 49476 2884 49478
rect 2778 48728 2834 48784
rect 2588 48442 2644 48444
rect 2668 48442 2724 48444
rect 2748 48442 2804 48444
rect 2828 48442 2884 48444
rect 2588 48390 2634 48442
rect 2634 48390 2644 48442
rect 2668 48390 2698 48442
rect 2698 48390 2710 48442
rect 2710 48390 2724 48442
rect 2748 48390 2762 48442
rect 2762 48390 2774 48442
rect 2774 48390 2804 48442
rect 2828 48390 2838 48442
rect 2838 48390 2884 48442
rect 2588 48388 2644 48390
rect 2668 48388 2724 48390
rect 2748 48388 2804 48390
rect 2828 48388 2884 48390
rect 2686 48220 2688 48240
rect 2688 48220 2740 48240
rect 2740 48220 2742 48240
rect 2686 48184 2742 48220
rect 3330 51176 3386 51232
rect 3054 50940 3056 50960
rect 3056 50940 3108 50960
rect 3108 50940 3110 50960
rect 3054 50904 3110 50940
rect 2588 47354 2644 47356
rect 2668 47354 2724 47356
rect 2748 47354 2804 47356
rect 2828 47354 2884 47356
rect 2588 47302 2634 47354
rect 2634 47302 2644 47354
rect 2668 47302 2698 47354
rect 2698 47302 2710 47354
rect 2710 47302 2724 47354
rect 2748 47302 2762 47354
rect 2762 47302 2774 47354
rect 2774 47302 2804 47354
rect 2828 47302 2838 47354
rect 2838 47302 2884 47354
rect 2588 47300 2644 47302
rect 2668 47300 2724 47302
rect 2748 47300 2804 47302
rect 2828 47300 2884 47302
rect 4219 74010 4275 74012
rect 4299 74010 4355 74012
rect 4379 74010 4435 74012
rect 4459 74010 4515 74012
rect 4219 73958 4265 74010
rect 4265 73958 4275 74010
rect 4299 73958 4329 74010
rect 4329 73958 4341 74010
rect 4341 73958 4355 74010
rect 4379 73958 4393 74010
rect 4393 73958 4405 74010
rect 4405 73958 4435 74010
rect 4459 73958 4469 74010
rect 4469 73958 4515 74010
rect 4219 73956 4275 73958
rect 4299 73956 4355 73958
rect 4379 73956 4435 73958
rect 4459 73956 4515 73958
rect 4219 72922 4275 72924
rect 4299 72922 4355 72924
rect 4379 72922 4435 72924
rect 4459 72922 4515 72924
rect 4219 72870 4265 72922
rect 4265 72870 4275 72922
rect 4299 72870 4329 72922
rect 4329 72870 4341 72922
rect 4341 72870 4355 72922
rect 4379 72870 4393 72922
rect 4393 72870 4405 72922
rect 4405 72870 4435 72922
rect 4459 72870 4469 72922
rect 4469 72870 4515 72922
rect 4219 72868 4275 72870
rect 4299 72868 4355 72870
rect 4379 72868 4435 72870
rect 4459 72868 4515 72870
rect 4219 71834 4275 71836
rect 4299 71834 4355 71836
rect 4379 71834 4435 71836
rect 4459 71834 4515 71836
rect 4219 71782 4265 71834
rect 4265 71782 4275 71834
rect 4299 71782 4329 71834
rect 4329 71782 4341 71834
rect 4341 71782 4355 71834
rect 4379 71782 4393 71834
rect 4393 71782 4405 71834
rect 4405 71782 4435 71834
rect 4459 71782 4469 71834
rect 4469 71782 4515 71834
rect 4219 71780 4275 71782
rect 4299 71780 4355 71782
rect 4379 71780 4435 71782
rect 4459 71780 4515 71782
rect 3974 69264 4030 69320
rect 3974 68448 4030 68504
rect 3330 50768 3386 50824
rect 3054 46688 3110 46744
rect 2588 46266 2644 46268
rect 2668 46266 2724 46268
rect 2748 46266 2804 46268
rect 2828 46266 2884 46268
rect 2588 46214 2634 46266
rect 2634 46214 2644 46266
rect 2668 46214 2698 46266
rect 2698 46214 2710 46266
rect 2710 46214 2724 46266
rect 2748 46214 2762 46266
rect 2762 46214 2774 46266
rect 2774 46214 2804 46266
rect 2828 46214 2838 46266
rect 2838 46214 2884 46266
rect 2588 46212 2644 46214
rect 2668 46212 2724 46214
rect 2748 46212 2804 46214
rect 2828 46212 2884 46214
rect 2962 45772 2964 45792
rect 2964 45772 3016 45792
rect 3016 45772 3018 45792
rect 2962 45736 3018 45772
rect 2588 45178 2644 45180
rect 2668 45178 2724 45180
rect 2748 45178 2804 45180
rect 2828 45178 2884 45180
rect 2588 45126 2634 45178
rect 2634 45126 2644 45178
rect 2668 45126 2698 45178
rect 2698 45126 2710 45178
rect 2710 45126 2724 45178
rect 2748 45126 2762 45178
rect 2762 45126 2774 45178
rect 2774 45126 2804 45178
rect 2828 45126 2838 45178
rect 2838 45126 2884 45178
rect 2588 45124 2644 45126
rect 2668 45124 2724 45126
rect 2748 45124 2804 45126
rect 2828 45124 2884 45126
rect 2588 44090 2644 44092
rect 2668 44090 2724 44092
rect 2748 44090 2804 44092
rect 2828 44090 2884 44092
rect 2588 44038 2634 44090
rect 2634 44038 2644 44090
rect 2668 44038 2698 44090
rect 2698 44038 2710 44090
rect 2710 44038 2724 44090
rect 2748 44038 2762 44090
rect 2762 44038 2774 44090
rect 2774 44038 2804 44090
rect 2828 44038 2838 44090
rect 2838 44038 2884 44090
rect 2588 44036 2644 44038
rect 2668 44036 2724 44038
rect 2748 44036 2804 44038
rect 2828 44036 2884 44038
rect 2870 43288 2926 43344
rect 2588 43002 2644 43004
rect 2668 43002 2724 43004
rect 2748 43002 2804 43004
rect 2828 43002 2884 43004
rect 2588 42950 2634 43002
rect 2634 42950 2644 43002
rect 2668 42950 2698 43002
rect 2698 42950 2710 43002
rect 2710 42950 2724 43002
rect 2748 42950 2762 43002
rect 2762 42950 2774 43002
rect 2774 42950 2804 43002
rect 2828 42950 2838 43002
rect 2838 42950 2884 43002
rect 2588 42948 2644 42950
rect 2668 42948 2724 42950
rect 2748 42948 2804 42950
rect 2828 42948 2884 42950
rect 2588 41914 2644 41916
rect 2668 41914 2724 41916
rect 2748 41914 2804 41916
rect 2828 41914 2884 41916
rect 2588 41862 2634 41914
rect 2634 41862 2644 41914
rect 2668 41862 2698 41914
rect 2698 41862 2710 41914
rect 2710 41862 2724 41914
rect 2748 41862 2762 41914
rect 2762 41862 2774 41914
rect 2774 41862 2804 41914
rect 2828 41862 2838 41914
rect 2838 41862 2884 41914
rect 2588 41860 2644 41862
rect 2668 41860 2724 41862
rect 2748 41860 2804 41862
rect 2828 41860 2884 41862
rect 2226 38392 2282 38448
rect 2410 38664 2466 38720
rect 2318 37576 2374 37632
rect 2226 36216 2282 36272
rect 2410 35808 2466 35864
rect 2318 33632 2374 33688
rect 2588 40826 2644 40828
rect 2668 40826 2724 40828
rect 2748 40826 2804 40828
rect 2828 40826 2884 40828
rect 2588 40774 2634 40826
rect 2634 40774 2644 40826
rect 2668 40774 2698 40826
rect 2698 40774 2710 40826
rect 2710 40774 2724 40826
rect 2748 40774 2762 40826
rect 2762 40774 2774 40826
rect 2774 40774 2804 40826
rect 2828 40774 2838 40826
rect 2838 40774 2884 40826
rect 2588 40772 2644 40774
rect 2668 40772 2724 40774
rect 2748 40772 2804 40774
rect 2828 40772 2884 40774
rect 2588 39738 2644 39740
rect 2668 39738 2724 39740
rect 2748 39738 2804 39740
rect 2828 39738 2884 39740
rect 2588 39686 2634 39738
rect 2634 39686 2644 39738
rect 2668 39686 2698 39738
rect 2698 39686 2710 39738
rect 2710 39686 2724 39738
rect 2748 39686 2762 39738
rect 2762 39686 2774 39738
rect 2774 39686 2804 39738
rect 2828 39686 2838 39738
rect 2838 39686 2884 39738
rect 2588 39684 2644 39686
rect 2668 39684 2724 39686
rect 2748 39684 2804 39686
rect 2828 39684 2884 39686
rect 3054 43596 3056 43616
rect 3056 43596 3108 43616
rect 3108 43596 3110 43616
rect 3054 43560 3110 43596
rect 3054 43288 3110 43344
rect 3054 40160 3110 40216
rect 2962 38800 3018 38856
rect 2962 38664 3018 38720
rect 2588 38650 2644 38652
rect 2668 38650 2724 38652
rect 2748 38650 2804 38652
rect 2828 38650 2884 38652
rect 2588 38598 2634 38650
rect 2634 38598 2644 38650
rect 2668 38598 2698 38650
rect 2698 38598 2710 38650
rect 2710 38598 2724 38650
rect 2748 38598 2762 38650
rect 2762 38598 2774 38650
rect 2774 38598 2804 38650
rect 2828 38598 2838 38650
rect 2838 38598 2884 38650
rect 2588 38596 2644 38598
rect 2668 38596 2724 38598
rect 2748 38596 2804 38598
rect 2828 38596 2884 38598
rect 2588 37562 2644 37564
rect 2668 37562 2724 37564
rect 2748 37562 2804 37564
rect 2828 37562 2884 37564
rect 2588 37510 2634 37562
rect 2634 37510 2644 37562
rect 2668 37510 2698 37562
rect 2698 37510 2710 37562
rect 2710 37510 2724 37562
rect 2748 37510 2762 37562
rect 2762 37510 2774 37562
rect 2774 37510 2804 37562
rect 2828 37510 2838 37562
rect 2838 37510 2884 37562
rect 2588 37508 2644 37510
rect 2668 37508 2724 37510
rect 2748 37508 2804 37510
rect 2828 37508 2884 37510
rect 2962 37168 3018 37224
rect 2588 36474 2644 36476
rect 2668 36474 2724 36476
rect 2748 36474 2804 36476
rect 2828 36474 2884 36476
rect 2588 36422 2634 36474
rect 2634 36422 2644 36474
rect 2668 36422 2698 36474
rect 2698 36422 2710 36474
rect 2710 36422 2724 36474
rect 2748 36422 2762 36474
rect 2762 36422 2774 36474
rect 2774 36422 2804 36474
rect 2828 36422 2838 36474
rect 2838 36422 2884 36474
rect 2588 36420 2644 36422
rect 2668 36420 2724 36422
rect 2748 36420 2804 36422
rect 2828 36420 2884 36422
rect 2588 35386 2644 35388
rect 2668 35386 2724 35388
rect 2748 35386 2804 35388
rect 2828 35386 2884 35388
rect 2588 35334 2634 35386
rect 2634 35334 2644 35386
rect 2668 35334 2698 35386
rect 2698 35334 2710 35386
rect 2710 35334 2724 35386
rect 2748 35334 2762 35386
rect 2762 35334 2774 35386
rect 2774 35334 2804 35386
rect 2828 35334 2838 35386
rect 2838 35334 2884 35386
rect 2588 35332 2644 35334
rect 2668 35332 2724 35334
rect 2748 35332 2804 35334
rect 2828 35332 2884 35334
rect 2588 34298 2644 34300
rect 2668 34298 2724 34300
rect 2748 34298 2804 34300
rect 2828 34298 2884 34300
rect 2588 34246 2634 34298
rect 2634 34246 2644 34298
rect 2668 34246 2698 34298
rect 2698 34246 2710 34298
rect 2710 34246 2724 34298
rect 2748 34246 2762 34298
rect 2762 34246 2774 34298
rect 2774 34246 2804 34298
rect 2828 34246 2838 34298
rect 2838 34246 2884 34298
rect 2588 34244 2644 34246
rect 2668 34244 2724 34246
rect 2748 34244 2804 34246
rect 2828 34244 2884 34246
rect 1398 25880 1454 25936
rect 1490 25472 1546 25528
rect 1490 23296 1546 23352
rect 1398 22888 1454 22944
rect 1766 29144 1822 29200
rect 2588 33210 2644 33212
rect 2668 33210 2724 33212
rect 2748 33210 2804 33212
rect 2828 33210 2884 33212
rect 2588 33158 2634 33210
rect 2634 33158 2644 33210
rect 2668 33158 2698 33210
rect 2698 33158 2710 33210
rect 2710 33158 2724 33210
rect 2748 33158 2762 33210
rect 2762 33158 2774 33210
rect 2774 33158 2804 33210
rect 2828 33158 2838 33210
rect 2838 33158 2884 33210
rect 2588 33156 2644 33158
rect 2668 33156 2724 33158
rect 2748 33156 2804 33158
rect 2828 33156 2884 33158
rect 3054 36644 3110 36680
rect 3054 36624 3056 36644
rect 3056 36624 3108 36644
rect 3108 36624 3110 36644
rect 3054 34448 3110 34504
rect 2318 32816 2374 32872
rect 2318 32544 2374 32600
rect 2502 32408 2558 32464
rect 2226 31728 2282 31784
rect 2226 31592 2282 31648
rect 2134 29280 2190 29336
rect 1398 17720 1454 17776
rect 2410 31456 2466 31512
rect 2410 31084 2412 31104
rect 2412 31084 2464 31104
rect 2464 31084 2466 31104
rect 2410 31048 2466 31084
rect 2318 30232 2374 30288
rect 2588 32122 2644 32124
rect 2668 32122 2724 32124
rect 2748 32122 2804 32124
rect 2828 32122 2884 32124
rect 2588 32070 2634 32122
rect 2634 32070 2644 32122
rect 2668 32070 2698 32122
rect 2698 32070 2710 32122
rect 2710 32070 2724 32122
rect 2748 32070 2762 32122
rect 2762 32070 2774 32122
rect 2774 32070 2804 32122
rect 2828 32070 2838 32122
rect 2838 32070 2884 32122
rect 2588 32068 2644 32070
rect 2668 32068 2724 32070
rect 2748 32068 2804 32070
rect 2828 32068 2884 32070
rect 2588 31034 2644 31036
rect 2668 31034 2724 31036
rect 2748 31034 2804 31036
rect 2828 31034 2884 31036
rect 2588 30982 2634 31034
rect 2634 30982 2644 31034
rect 2668 30982 2698 31034
rect 2698 30982 2710 31034
rect 2710 30982 2724 31034
rect 2748 30982 2762 31034
rect 2762 30982 2774 31034
rect 2774 30982 2804 31034
rect 2828 30982 2838 31034
rect 2838 30982 2884 31034
rect 2588 30980 2644 30982
rect 2668 30980 2724 30982
rect 2748 30980 2804 30982
rect 2828 30980 2884 30982
rect 2588 29946 2644 29948
rect 2668 29946 2724 29948
rect 2748 29946 2804 29948
rect 2828 29946 2884 29948
rect 2588 29894 2634 29946
rect 2634 29894 2644 29946
rect 2668 29894 2698 29946
rect 2698 29894 2710 29946
rect 2710 29894 2724 29946
rect 2748 29894 2762 29946
rect 2762 29894 2774 29946
rect 2774 29894 2804 29946
rect 2828 29894 2838 29946
rect 2838 29894 2884 29946
rect 2588 29892 2644 29894
rect 2668 29892 2724 29894
rect 2748 29892 2804 29894
rect 2828 29892 2884 29894
rect 2962 29688 3018 29744
rect 2778 28952 2834 29008
rect 2588 28858 2644 28860
rect 2668 28858 2724 28860
rect 2748 28858 2804 28860
rect 2828 28858 2884 28860
rect 2588 28806 2634 28858
rect 2634 28806 2644 28858
rect 2668 28806 2698 28858
rect 2698 28806 2710 28858
rect 2710 28806 2724 28858
rect 2748 28806 2762 28858
rect 2762 28806 2774 28858
rect 2774 28806 2804 28858
rect 2828 28806 2838 28858
rect 2838 28806 2884 28858
rect 2588 28804 2644 28806
rect 2668 28804 2724 28806
rect 2748 28804 2804 28806
rect 2828 28804 2884 28806
rect 2134 25880 2190 25936
rect 1398 12280 1454 12336
rect 1490 11736 1546 11792
rect 1398 11328 1454 11384
rect 1306 10920 1362 10976
rect 1398 10376 1454 10432
rect 1306 9968 1362 10024
rect 1398 9560 1454 9616
rect 1398 9152 1454 9208
rect 1858 15136 1914 15192
rect 2588 27770 2644 27772
rect 2668 27770 2724 27772
rect 2748 27770 2804 27772
rect 2828 27770 2884 27772
rect 2588 27718 2634 27770
rect 2634 27718 2644 27770
rect 2668 27718 2698 27770
rect 2698 27718 2710 27770
rect 2710 27718 2724 27770
rect 2748 27718 2762 27770
rect 2762 27718 2774 27770
rect 2774 27718 2804 27770
rect 2828 27718 2838 27770
rect 2838 27718 2884 27770
rect 2588 27716 2644 27718
rect 2668 27716 2724 27718
rect 2748 27716 2804 27718
rect 2828 27716 2884 27718
rect 2778 27512 2834 27568
rect 2870 27376 2926 27432
rect 2588 26682 2644 26684
rect 2668 26682 2724 26684
rect 2748 26682 2804 26684
rect 2828 26682 2884 26684
rect 2588 26630 2634 26682
rect 2634 26630 2644 26682
rect 2668 26630 2698 26682
rect 2698 26630 2710 26682
rect 2710 26630 2724 26682
rect 2748 26630 2762 26682
rect 2762 26630 2774 26682
rect 2774 26630 2804 26682
rect 2828 26630 2838 26682
rect 2838 26630 2884 26682
rect 2588 26628 2644 26630
rect 2668 26628 2724 26630
rect 2748 26628 2804 26630
rect 2828 26628 2884 26630
rect 2588 25594 2644 25596
rect 2668 25594 2724 25596
rect 2748 25594 2804 25596
rect 2828 25594 2884 25596
rect 2588 25542 2634 25594
rect 2634 25542 2644 25594
rect 2668 25542 2698 25594
rect 2698 25542 2710 25594
rect 2710 25542 2724 25594
rect 2748 25542 2762 25594
rect 2762 25542 2774 25594
rect 2774 25542 2804 25594
rect 2828 25542 2838 25594
rect 2838 25542 2884 25594
rect 2588 25540 2644 25542
rect 2668 25540 2724 25542
rect 2748 25540 2804 25542
rect 2828 25540 2884 25542
rect 2594 25336 2650 25392
rect 2962 25064 3018 25120
rect 2588 24506 2644 24508
rect 2668 24506 2724 24508
rect 2748 24506 2804 24508
rect 2828 24506 2884 24508
rect 2588 24454 2634 24506
rect 2634 24454 2644 24506
rect 2668 24454 2698 24506
rect 2698 24454 2710 24506
rect 2710 24454 2724 24506
rect 2748 24454 2762 24506
rect 2762 24454 2774 24506
rect 2774 24454 2804 24506
rect 2828 24454 2838 24506
rect 2838 24454 2884 24506
rect 2588 24452 2644 24454
rect 2668 24452 2724 24454
rect 2748 24452 2804 24454
rect 2828 24452 2884 24454
rect 2588 23418 2644 23420
rect 2668 23418 2724 23420
rect 2748 23418 2804 23420
rect 2828 23418 2884 23420
rect 2588 23366 2634 23418
rect 2634 23366 2644 23418
rect 2668 23366 2698 23418
rect 2698 23366 2710 23418
rect 2710 23366 2724 23418
rect 2748 23366 2762 23418
rect 2762 23366 2774 23418
rect 2774 23366 2804 23418
rect 2828 23366 2838 23418
rect 2838 23366 2884 23418
rect 2588 23364 2644 23366
rect 2668 23364 2724 23366
rect 2748 23364 2804 23366
rect 2828 23364 2884 23366
rect 2588 22330 2644 22332
rect 2668 22330 2724 22332
rect 2748 22330 2804 22332
rect 2828 22330 2884 22332
rect 2588 22278 2634 22330
rect 2634 22278 2644 22330
rect 2668 22278 2698 22330
rect 2698 22278 2710 22330
rect 2710 22278 2724 22330
rect 2748 22278 2762 22330
rect 2762 22278 2774 22330
rect 2774 22278 2804 22330
rect 2828 22278 2838 22330
rect 2838 22278 2884 22330
rect 2588 22276 2644 22278
rect 2668 22276 2724 22278
rect 2748 22276 2804 22278
rect 2828 22276 2884 22278
rect 2870 21392 2926 21448
rect 2588 21242 2644 21244
rect 2668 21242 2724 21244
rect 2748 21242 2804 21244
rect 2828 21242 2884 21244
rect 2588 21190 2634 21242
rect 2634 21190 2644 21242
rect 2668 21190 2698 21242
rect 2698 21190 2710 21242
rect 2710 21190 2724 21242
rect 2748 21190 2762 21242
rect 2762 21190 2774 21242
rect 2774 21190 2804 21242
rect 2828 21190 2838 21242
rect 2838 21190 2884 21242
rect 2588 21188 2644 21190
rect 2668 21188 2724 21190
rect 2748 21188 2804 21190
rect 2828 21188 2884 21190
rect 2226 16496 2282 16552
rect 2588 20154 2644 20156
rect 2668 20154 2724 20156
rect 2748 20154 2804 20156
rect 2828 20154 2884 20156
rect 2588 20102 2634 20154
rect 2634 20102 2644 20154
rect 2668 20102 2698 20154
rect 2698 20102 2710 20154
rect 2710 20102 2724 20154
rect 2748 20102 2762 20154
rect 2762 20102 2774 20154
rect 2774 20102 2804 20154
rect 2828 20102 2838 20154
rect 2838 20102 2884 20154
rect 2588 20100 2644 20102
rect 2668 20100 2724 20102
rect 2748 20100 2804 20102
rect 2828 20100 2884 20102
rect 2588 19066 2644 19068
rect 2668 19066 2724 19068
rect 2748 19066 2804 19068
rect 2828 19066 2884 19068
rect 2588 19014 2634 19066
rect 2634 19014 2644 19066
rect 2668 19014 2698 19066
rect 2698 19014 2710 19066
rect 2710 19014 2724 19066
rect 2748 19014 2762 19066
rect 2762 19014 2774 19066
rect 2774 19014 2804 19066
rect 2828 19014 2838 19066
rect 2838 19014 2884 19066
rect 2588 19012 2644 19014
rect 2668 19012 2724 19014
rect 2748 19012 2804 19014
rect 2828 19012 2884 19014
rect 2778 18128 2834 18184
rect 2588 17978 2644 17980
rect 2668 17978 2724 17980
rect 2748 17978 2804 17980
rect 2828 17978 2884 17980
rect 2588 17926 2634 17978
rect 2634 17926 2644 17978
rect 2668 17926 2698 17978
rect 2698 17926 2710 17978
rect 2710 17926 2724 17978
rect 2748 17926 2762 17978
rect 2762 17926 2774 17978
rect 2774 17926 2804 17978
rect 2828 17926 2838 17978
rect 2838 17926 2884 17978
rect 2588 17924 2644 17926
rect 2668 17924 2724 17926
rect 2748 17924 2804 17926
rect 2828 17924 2884 17926
rect 3422 45600 3478 45656
rect 3238 34040 3294 34096
rect 3698 57568 3754 57624
rect 3882 63844 3938 63880
rect 3882 63824 3884 63844
rect 3884 63824 3936 63844
rect 3936 63824 3938 63844
rect 4219 70746 4275 70748
rect 4299 70746 4355 70748
rect 4379 70746 4435 70748
rect 4459 70746 4515 70748
rect 4219 70694 4265 70746
rect 4265 70694 4275 70746
rect 4299 70694 4329 70746
rect 4329 70694 4341 70746
rect 4341 70694 4355 70746
rect 4379 70694 4393 70746
rect 4393 70694 4405 70746
rect 4405 70694 4435 70746
rect 4459 70694 4469 70746
rect 4469 70694 4515 70746
rect 4219 70692 4275 70694
rect 4299 70692 4355 70694
rect 4379 70692 4435 70694
rect 4459 70692 4515 70694
rect 4219 69658 4275 69660
rect 4299 69658 4355 69660
rect 4379 69658 4435 69660
rect 4459 69658 4515 69660
rect 4219 69606 4265 69658
rect 4265 69606 4275 69658
rect 4299 69606 4329 69658
rect 4329 69606 4341 69658
rect 4341 69606 4355 69658
rect 4379 69606 4393 69658
rect 4393 69606 4405 69658
rect 4405 69606 4435 69658
rect 4459 69606 4469 69658
rect 4469 69606 4515 69658
rect 4219 69604 4275 69606
rect 4299 69604 4355 69606
rect 4379 69604 4435 69606
rect 4459 69604 4515 69606
rect 4158 68856 4214 68912
rect 4219 68570 4275 68572
rect 4299 68570 4355 68572
rect 4379 68570 4435 68572
rect 4459 68570 4515 68572
rect 4219 68518 4265 68570
rect 4265 68518 4275 68570
rect 4299 68518 4329 68570
rect 4329 68518 4341 68570
rect 4341 68518 4355 68570
rect 4379 68518 4393 68570
rect 4393 68518 4405 68570
rect 4405 68518 4435 68570
rect 4459 68518 4469 68570
rect 4469 68518 4515 68570
rect 4219 68516 4275 68518
rect 4299 68516 4355 68518
rect 4379 68516 4435 68518
rect 4459 68516 4515 68518
rect 4219 67482 4275 67484
rect 4299 67482 4355 67484
rect 4379 67482 4435 67484
rect 4459 67482 4515 67484
rect 4219 67430 4265 67482
rect 4265 67430 4275 67482
rect 4299 67430 4329 67482
rect 4329 67430 4341 67482
rect 4341 67430 4355 67482
rect 4379 67430 4393 67482
rect 4393 67430 4405 67482
rect 4405 67430 4435 67482
rect 4459 67430 4469 67482
rect 4469 67430 4515 67482
rect 4219 67428 4275 67430
rect 4299 67428 4355 67430
rect 4379 67428 4435 67430
rect 4459 67428 4515 67430
rect 4219 66394 4275 66396
rect 4299 66394 4355 66396
rect 4379 66394 4435 66396
rect 4459 66394 4515 66396
rect 4219 66342 4265 66394
rect 4265 66342 4275 66394
rect 4299 66342 4329 66394
rect 4329 66342 4341 66394
rect 4341 66342 4355 66394
rect 4379 66342 4393 66394
rect 4393 66342 4405 66394
rect 4405 66342 4435 66394
rect 4459 66342 4469 66394
rect 4469 66342 4515 66394
rect 4219 66340 4275 66342
rect 4299 66340 4355 66342
rect 4379 66340 4435 66342
rect 4459 66340 4515 66342
rect 4219 65306 4275 65308
rect 4299 65306 4355 65308
rect 4379 65306 4435 65308
rect 4459 65306 4515 65308
rect 4219 65254 4265 65306
rect 4265 65254 4275 65306
rect 4299 65254 4329 65306
rect 4329 65254 4341 65306
rect 4341 65254 4355 65306
rect 4379 65254 4393 65306
rect 4393 65254 4405 65306
rect 4405 65254 4435 65306
rect 4459 65254 4469 65306
rect 4469 65254 4515 65306
rect 4219 65252 4275 65254
rect 4299 65252 4355 65254
rect 4379 65252 4435 65254
rect 4459 65252 4515 65254
rect 4219 64218 4275 64220
rect 4299 64218 4355 64220
rect 4379 64218 4435 64220
rect 4459 64218 4515 64220
rect 4219 64166 4265 64218
rect 4265 64166 4275 64218
rect 4299 64166 4329 64218
rect 4329 64166 4341 64218
rect 4341 64166 4355 64218
rect 4379 64166 4393 64218
rect 4393 64166 4405 64218
rect 4405 64166 4435 64218
rect 4459 64166 4469 64218
rect 4469 64166 4515 64218
rect 4219 64164 4275 64166
rect 4299 64164 4355 64166
rect 4379 64164 4435 64166
rect 4459 64164 4515 64166
rect 4066 63416 4122 63472
rect 4066 63144 4122 63200
rect 4219 63130 4275 63132
rect 4299 63130 4355 63132
rect 4379 63130 4435 63132
rect 4459 63130 4515 63132
rect 4219 63078 4265 63130
rect 4265 63078 4275 63130
rect 4299 63078 4329 63130
rect 4329 63078 4341 63130
rect 4341 63078 4355 63130
rect 4379 63078 4393 63130
rect 4393 63078 4405 63130
rect 4405 63078 4435 63130
rect 4459 63078 4469 63130
rect 4469 63078 4515 63130
rect 4219 63076 4275 63078
rect 4299 63076 4355 63078
rect 4379 63076 4435 63078
rect 4459 63076 4515 63078
rect 3974 62872 4030 62928
rect 4219 62042 4275 62044
rect 4299 62042 4355 62044
rect 4379 62042 4435 62044
rect 4459 62042 4515 62044
rect 4219 61990 4265 62042
rect 4265 61990 4275 62042
rect 4299 61990 4329 62042
rect 4329 61990 4341 62042
rect 4341 61990 4355 62042
rect 4379 61990 4393 62042
rect 4393 61990 4405 62042
rect 4405 61990 4435 62042
rect 4459 61990 4469 62042
rect 4469 61990 4515 62042
rect 4219 61988 4275 61990
rect 4299 61988 4355 61990
rect 4379 61988 4435 61990
rect 4459 61988 4515 61990
rect 3974 61104 4030 61160
rect 3882 60696 3938 60752
rect 3974 55564 3976 55584
rect 3976 55564 4028 55584
rect 4028 55564 4030 55584
rect 3974 55528 4030 55564
rect 3698 51060 3754 51096
rect 3698 51040 3700 51060
rect 3700 51040 3752 51060
rect 3752 51040 3754 51060
rect 3790 50496 3846 50552
rect 3882 49544 3938 49600
rect 3882 49136 3938 49192
rect 3790 44920 3846 44976
rect 3606 44376 3662 44432
rect 3514 39888 3570 39944
rect 4219 60954 4275 60956
rect 4299 60954 4355 60956
rect 4379 60954 4435 60956
rect 4459 60954 4515 60956
rect 4219 60902 4265 60954
rect 4265 60902 4275 60954
rect 4299 60902 4329 60954
rect 4329 60902 4341 60954
rect 4341 60902 4355 60954
rect 4379 60902 4393 60954
rect 4393 60902 4405 60954
rect 4405 60902 4435 60954
rect 4459 60902 4469 60954
rect 4469 60902 4515 60954
rect 4219 60900 4275 60902
rect 4299 60900 4355 60902
rect 4379 60900 4435 60902
rect 4459 60900 4515 60902
rect 4219 59866 4275 59868
rect 4299 59866 4355 59868
rect 4379 59866 4435 59868
rect 4459 59866 4515 59868
rect 4219 59814 4265 59866
rect 4265 59814 4275 59866
rect 4299 59814 4329 59866
rect 4329 59814 4341 59866
rect 4341 59814 4355 59866
rect 4379 59814 4393 59866
rect 4393 59814 4405 59866
rect 4405 59814 4435 59866
rect 4459 59814 4469 59866
rect 4469 59814 4515 59866
rect 4219 59812 4275 59814
rect 4299 59812 4355 59814
rect 4379 59812 4435 59814
rect 4459 59812 4515 59814
rect 4219 58778 4275 58780
rect 4299 58778 4355 58780
rect 4379 58778 4435 58780
rect 4459 58778 4515 58780
rect 4219 58726 4265 58778
rect 4265 58726 4275 58778
rect 4299 58726 4329 58778
rect 4329 58726 4341 58778
rect 4341 58726 4355 58778
rect 4379 58726 4393 58778
rect 4393 58726 4405 58778
rect 4405 58726 4435 58778
rect 4459 58726 4469 58778
rect 4469 58726 4515 58778
rect 4219 58724 4275 58726
rect 4299 58724 4355 58726
rect 4379 58724 4435 58726
rect 4459 58724 4515 58726
rect 4219 57690 4275 57692
rect 4299 57690 4355 57692
rect 4379 57690 4435 57692
rect 4459 57690 4515 57692
rect 4219 57638 4265 57690
rect 4265 57638 4275 57690
rect 4299 57638 4329 57690
rect 4329 57638 4341 57690
rect 4341 57638 4355 57690
rect 4379 57638 4393 57690
rect 4393 57638 4405 57690
rect 4405 57638 4435 57690
rect 4459 57638 4469 57690
rect 4469 57638 4515 57690
rect 4219 57636 4275 57638
rect 4299 57636 4355 57638
rect 4379 57636 4435 57638
rect 4459 57636 4515 57638
rect 4219 56602 4275 56604
rect 4299 56602 4355 56604
rect 4379 56602 4435 56604
rect 4459 56602 4515 56604
rect 4219 56550 4265 56602
rect 4265 56550 4275 56602
rect 4299 56550 4329 56602
rect 4329 56550 4341 56602
rect 4341 56550 4355 56602
rect 4379 56550 4393 56602
rect 4393 56550 4405 56602
rect 4405 56550 4435 56602
rect 4459 56550 4469 56602
rect 4469 56550 4515 56602
rect 4219 56548 4275 56550
rect 4299 56548 4355 56550
rect 4379 56548 4435 56550
rect 4459 56548 4515 56550
rect 4219 55514 4275 55516
rect 4299 55514 4355 55516
rect 4379 55514 4435 55516
rect 4459 55514 4515 55516
rect 4219 55462 4265 55514
rect 4265 55462 4275 55514
rect 4299 55462 4329 55514
rect 4329 55462 4341 55514
rect 4341 55462 4355 55514
rect 4379 55462 4393 55514
rect 4393 55462 4405 55514
rect 4405 55462 4435 55514
rect 4459 55462 4469 55514
rect 4469 55462 4515 55514
rect 4219 55460 4275 55462
rect 4299 55460 4355 55462
rect 4379 55460 4435 55462
rect 4459 55460 4515 55462
rect 4219 54426 4275 54428
rect 4299 54426 4355 54428
rect 4379 54426 4435 54428
rect 4459 54426 4515 54428
rect 4219 54374 4265 54426
rect 4265 54374 4275 54426
rect 4299 54374 4329 54426
rect 4329 54374 4341 54426
rect 4341 54374 4355 54426
rect 4379 54374 4393 54426
rect 4393 54374 4405 54426
rect 4405 54374 4435 54426
rect 4459 54374 4469 54426
rect 4469 54374 4515 54426
rect 4219 54372 4275 54374
rect 4299 54372 4355 54374
rect 4379 54372 4435 54374
rect 4459 54372 4515 54374
rect 4219 53338 4275 53340
rect 4299 53338 4355 53340
rect 4379 53338 4435 53340
rect 4459 53338 4515 53340
rect 4219 53286 4265 53338
rect 4265 53286 4275 53338
rect 4299 53286 4329 53338
rect 4329 53286 4341 53338
rect 4341 53286 4355 53338
rect 4379 53286 4393 53338
rect 4393 53286 4405 53338
rect 4405 53286 4435 53338
rect 4459 53286 4469 53338
rect 4469 53286 4515 53338
rect 4219 53284 4275 53286
rect 4299 53284 4355 53286
rect 4379 53284 4435 53286
rect 4459 53284 4515 53286
rect 4219 52250 4275 52252
rect 4299 52250 4355 52252
rect 4379 52250 4435 52252
rect 4459 52250 4515 52252
rect 4219 52198 4265 52250
rect 4265 52198 4275 52250
rect 4299 52198 4329 52250
rect 4329 52198 4341 52250
rect 4341 52198 4355 52250
rect 4379 52198 4393 52250
rect 4393 52198 4405 52250
rect 4405 52198 4435 52250
rect 4459 52198 4469 52250
rect 4469 52198 4515 52250
rect 4219 52196 4275 52198
rect 4299 52196 4355 52198
rect 4379 52196 4435 52198
rect 4459 52196 4515 52198
rect 4219 51162 4275 51164
rect 4299 51162 4355 51164
rect 4379 51162 4435 51164
rect 4459 51162 4515 51164
rect 4219 51110 4265 51162
rect 4265 51110 4275 51162
rect 4299 51110 4329 51162
rect 4329 51110 4341 51162
rect 4341 51110 4355 51162
rect 4379 51110 4393 51162
rect 4393 51110 4405 51162
rect 4405 51110 4435 51162
rect 4459 51110 4469 51162
rect 4469 51110 4515 51162
rect 4219 51108 4275 51110
rect 4299 51108 4355 51110
rect 4379 51108 4435 51110
rect 4459 51108 4515 51110
rect 4219 50074 4275 50076
rect 4299 50074 4355 50076
rect 4379 50074 4435 50076
rect 4459 50074 4515 50076
rect 4219 50022 4265 50074
rect 4265 50022 4275 50074
rect 4299 50022 4329 50074
rect 4329 50022 4341 50074
rect 4341 50022 4355 50074
rect 4379 50022 4393 50074
rect 4393 50022 4405 50074
rect 4405 50022 4435 50074
rect 4459 50022 4469 50074
rect 4469 50022 4515 50074
rect 4219 50020 4275 50022
rect 4299 50020 4355 50022
rect 4379 50020 4435 50022
rect 4459 50020 4515 50022
rect 4158 49852 4160 49872
rect 4160 49852 4212 49872
rect 4212 49852 4214 49872
rect 4158 49816 4214 49852
rect 4219 48986 4275 48988
rect 4299 48986 4355 48988
rect 4379 48986 4435 48988
rect 4459 48986 4515 48988
rect 4219 48934 4265 48986
rect 4265 48934 4275 48986
rect 4299 48934 4329 48986
rect 4329 48934 4341 48986
rect 4341 48934 4355 48986
rect 4379 48934 4393 48986
rect 4393 48934 4405 48986
rect 4405 48934 4435 48986
rect 4459 48934 4469 48986
rect 4469 48934 4515 48986
rect 4219 48932 4275 48934
rect 4299 48932 4355 48934
rect 4379 48932 4435 48934
rect 4459 48932 4515 48934
rect 5851 74554 5907 74556
rect 5931 74554 5987 74556
rect 6011 74554 6067 74556
rect 6091 74554 6147 74556
rect 5851 74502 5897 74554
rect 5897 74502 5907 74554
rect 5931 74502 5961 74554
rect 5961 74502 5973 74554
rect 5973 74502 5987 74554
rect 6011 74502 6025 74554
rect 6025 74502 6037 74554
rect 6037 74502 6067 74554
rect 6091 74502 6101 74554
rect 6101 74502 6147 74554
rect 5851 74500 5907 74502
rect 5931 74500 5987 74502
rect 6011 74500 6067 74502
rect 6091 74500 6147 74502
rect 4219 47898 4275 47900
rect 4299 47898 4355 47900
rect 4379 47898 4435 47900
rect 4459 47898 4515 47900
rect 4219 47846 4265 47898
rect 4265 47846 4275 47898
rect 4299 47846 4329 47898
rect 4329 47846 4341 47898
rect 4341 47846 4355 47898
rect 4379 47846 4393 47898
rect 4393 47846 4405 47898
rect 4405 47846 4435 47898
rect 4459 47846 4469 47898
rect 4469 47846 4515 47898
rect 4219 47844 4275 47846
rect 4299 47844 4355 47846
rect 4379 47844 4435 47846
rect 4459 47844 4515 47846
rect 4219 46810 4275 46812
rect 4299 46810 4355 46812
rect 4379 46810 4435 46812
rect 4459 46810 4515 46812
rect 4219 46758 4265 46810
rect 4265 46758 4275 46810
rect 4299 46758 4329 46810
rect 4329 46758 4341 46810
rect 4341 46758 4355 46810
rect 4379 46758 4393 46810
rect 4393 46758 4405 46810
rect 4405 46758 4435 46810
rect 4459 46758 4469 46810
rect 4469 46758 4515 46810
rect 4219 46756 4275 46758
rect 4299 46756 4355 46758
rect 4379 46756 4435 46758
rect 4459 46756 4515 46758
rect 4802 49544 4858 49600
rect 4219 45722 4275 45724
rect 4299 45722 4355 45724
rect 4379 45722 4435 45724
rect 4459 45722 4515 45724
rect 4219 45670 4265 45722
rect 4265 45670 4275 45722
rect 4299 45670 4329 45722
rect 4329 45670 4341 45722
rect 4341 45670 4355 45722
rect 4379 45670 4393 45722
rect 4393 45670 4405 45722
rect 4405 45670 4435 45722
rect 4459 45670 4469 45722
rect 4469 45670 4515 45722
rect 4219 45668 4275 45670
rect 4299 45668 4355 45670
rect 4379 45668 4435 45670
rect 4459 45668 4515 45670
rect 4219 44634 4275 44636
rect 4299 44634 4355 44636
rect 4379 44634 4435 44636
rect 4459 44634 4515 44636
rect 4219 44582 4265 44634
rect 4265 44582 4275 44634
rect 4299 44582 4329 44634
rect 4329 44582 4341 44634
rect 4341 44582 4355 44634
rect 4379 44582 4393 44634
rect 4393 44582 4405 44634
rect 4405 44582 4435 44634
rect 4459 44582 4469 44634
rect 4469 44582 4515 44634
rect 4219 44580 4275 44582
rect 4299 44580 4355 44582
rect 4379 44580 4435 44582
rect 4459 44580 4515 44582
rect 4219 43546 4275 43548
rect 4299 43546 4355 43548
rect 4379 43546 4435 43548
rect 4459 43546 4515 43548
rect 4219 43494 4265 43546
rect 4265 43494 4275 43546
rect 4299 43494 4329 43546
rect 4329 43494 4341 43546
rect 4341 43494 4355 43546
rect 4379 43494 4393 43546
rect 4393 43494 4405 43546
rect 4405 43494 4435 43546
rect 4459 43494 4469 43546
rect 4469 43494 4515 43546
rect 4219 43492 4275 43494
rect 4299 43492 4355 43494
rect 4379 43492 4435 43494
rect 4459 43492 4515 43494
rect 4526 43288 4582 43344
rect 4219 42458 4275 42460
rect 4299 42458 4355 42460
rect 4379 42458 4435 42460
rect 4459 42458 4515 42460
rect 4219 42406 4265 42458
rect 4265 42406 4275 42458
rect 4299 42406 4329 42458
rect 4329 42406 4341 42458
rect 4341 42406 4355 42458
rect 4379 42406 4393 42458
rect 4393 42406 4405 42458
rect 4405 42406 4435 42458
rect 4459 42406 4469 42458
rect 4469 42406 4515 42458
rect 4219 42404 4275 42406
rect 4299 42404 4355 42406
rect 4379 42404 4435 42406
rect 4459 42404 4515 42406
rect 4158 42200 4214 42256
rect 4219 41370 4275 41372
rect 4299 41370 4355 41372
rect 4379 41370 4435 41372
rect 4459 41370 4515 41372
rect 4219 41318 4265 41370
rect 4265 41318 4275 41370
rect 4299 41318 4329 41370
rect 4329 41318 4341 41370
rect 4341 41318 4355 41370
rect 4379 41318 4393 41370
rect 4393 41318 4405 41370
rect 4405 41318 4435 41370
rect 4459 41318 4469 41370
rect 4469 41318 4515 41370
rect 4219 41316 4275 41318
rect 4299 41316 4355 41318
rect 4379 41316 4435 41318
rect 4459 41316 4515 41318
rect 4219 40282 4275 40284
rect 4299 40282 4355 40284
rect 4379 40282 4435 40284
rect 4459 40282 4515 40284
rect 4219 40230 4265 40282
rect 4265 40230 4275 40282
rect 4299 40230 4329 40282
rect 4329 40230 4341 40282
rect 4341 40230 4355 40282
rect 4379 40230 4393 40282
rect 4393 40230 4405 40282
rect 4405 40230 4435 40282
rect 4459 40230 4469 40282
rect 4469 40230 4515 40282
rect 4219 40228 4275 40230
rect 4299 40228 4355 40230
rect 4379 40228 4435 40230
rect 4459 40228 4515 40230
rect 3882 39480 3938 39536
rect 3514 36896 3570 36952
rect 3514 36624 3570 36680
rect 3330 33768 3386 33824
rect 3422 28464 3478 28520
rect 3422 27240 3478 27296
rect 4066 40024 4122 40080
rect 4219 39194 4275 39196
rect 4299 39194 4355 39196
rect 4379 39194 4435 39196
rect 4459 39194 4515 39196
rect 4219 39142 4265 39194
rect 4265 39142 4275 39194
rect 4299 39142 4329 39194
rect 4329 39142 4341 39194
rect 4341 39142 4355 39194
rect 4379 39142 4393 39194
rect 4393 39142 4405 39194
rect 4405 39142 4435 39194
rect 4459 39142 4469 39194
rect 4469 39142 4515 39194
rect 4219 39140 4275 39142
rect 4299 39140 4355 39142
rect 4379 39140 4435 39142
rect 4459 39140 4515 39142
rect 4066 38956 4122 38992
rect 4066 38936 4068 38956
rect 4068 38936 4120 38956
rect 4120 38936 4122 38956
rect 4342 38800 4398 38856
rect 3974 37304 4030 37360
rect 3882 36896 3938 36952
rect 3698 35400 3754 35456
rect 3606 31592 3662 31648
rect 4219 38106 4275 38108
rect 4299 38106 4355 38108
rect 4379 38106 4435 38108
rect 4459 38106 4515 38108
rect 4219 38054 4265 38106
rect 4265 38054 4275 38106
rect 4299 38054 4329 38106
rect 4329 38054 4341 38106
rect 4341 38054 4355 38106
rect 4379 38054 4393 38106
rect 4393 38054 4405 38106
rect 4405 38054 4435 38106
rect 4459 38054 4469 38106
rect 4469 38054 4515 38106
rect 4219 38052 4275 38054
rect 4299 38052 4355 38054
rect 4379 38052 4435 38054
rect 4459 38052 4515 38054
rect 4219 37018 4275 37020
rect 4299 37018 4355 37020
rect 4379 37018 4435 37020
rect 4459 37018 4515 37020
rect 4219 36966 4265 37018
rect 4265 36966 4275 37018
rect 4299 36966 4329 37018
rect 4329 36966 4341 37018
rect 4341 36966 4355 37018
rect 4379 36966 4393 37018
rect 4393 36966 4405 37018
rect 4405 36966 4435 37018
rect 4459 36966 4469 37018
rect 4469 36966 4515 37018
rect 4219 36964 4275 36966
rect 4299 36964 4355 36966
rect 4379 36964 4435 36966
rect 4459 36964 4515 36966
rect 3790 28600 3846 28656
rect 3698 26868 3700 26888
rect 3700 26868 3752 26888
rect 3752 26868 3754 26888
rect 3238 24656 3294 24712
rect 3146 23704 3202 23760
rect 3146 22480 3202 22536
rect 3698 26832 3754 26868
rect 3606 26732 3608 26752
rect 3608 26732 3660 26752
rect 3660 26732 3662 26752
rect 3606 26696 3662 26732
rect 3514 26324 3516 26344
rect 3516 26324 3568 26344
rect 3568 26324 3570 26344
rect 3514 26288 3570 26324
rect 3054 19216 3110 19272
rect 3238 18536 3294 18592
rect 2870 17040 2926 17096
rect 2588 16890 2644 16892
rect 2668 16890 2724 16892
rect 2748 16890 2804 16892
rect 2828 16890 2884 16892
rect 2588 16838 2634 16890
rect 2634 16838 2644 16890
rect 2668 16838 2698 16890
rect 2698 16838 2710 16890
rect 2710 16838 2724 16890
rect 2748 16838 2762 16890
rect 2762 16838 2774 16890
rect 2774 16838 2804 16890
rect 2828 16838 2838 16890
rect 2838 16838 2884 16890
rect 2588 16836 2644 16838
rect 2668 16836 2724 16838
rect 2748 16836 2804 16838
rect 2828 16836 2884 16838
rect 3054 17312 3110 17368
rect 2588 15802 2644 15804
rect 2668 15802 2724 15804
rect 2748 15802 2804 15804
rect 2828 15802 2884 15804
rect 2588 15750 2634 15802
rect 2634 15750 2644 15802
rect 2668 15750 2698 15802
rect 2698 15750 2710 15802
rect 2710 15750 2724 15802
rect 2748 15750 2762 15802
rect 2762 15750 2774 15802
rect 2774 15750 2804 15802
rect 2828 15750 2838 15802
rect 2838 15750 2884 15802
rect 2588 15748 2644 15750
rect 2668 15748 2724 15750
rect 2748 15748 2804 15750
rect 2828 15748 2884 15750
rect 1858 12960 1914 13016
rect 1398 8336 1454 8392
rect 1306 7792 1362 7848
rect 1398 7384 1454 7440
rect 1858 6568 1914 6624
rect 1306 3168 1362 3224
rect 1398 2624 1454 2680
rect 2778 15156 2834 15192
rect 2778 15136 2780 15156
rect 2780 15136 2832 15156
rect 2832 15136 2834 15156
rect 2588 14714 2644 14716
rect 2668 14714 2724 14716
rect 2748 14714 2804 14716
rect 2828 14714 2884 14716
rect 2588 14662 2634 14714
rect 2634 14662 2644 14714
rect 2668 14662 2698 14714
rect 2698 14662 2710 14714
rect 2710 14662 2724 14714
rect 2748 14662 2762 14714
rect 2762 14662 2774 14714
rect 2774 14662 2804 14714
rect 2828 14662 2838 14714
rect 2838 14662 2884 14714
rect 2588 14660 2644 14662
rect 2668 14660 2724 14662
rect 2748 14660 2804 14662
rect 2828 14660 2884 14662
rect 2588 13626 2644 13628
rect 2668 13626 2724 13628
rect 2748 13626 2804 13628
rect 2828 13626 2884 13628
rect 2588 13574 2634 13626
rect 2634 13574 2644 13626
rect 2668 13574 2698 13626
rect 2698 13574 2710 13626
rect 2710 13574 2724 13626
rect 2748 13574 2762 13626
rect 2762 13574 2774 13626
rect 2774 13574 2804 13626
rect 2828 13574 2838 13626
rect 2838 13574 2884 13626
rect 2588 13572 2644 13574
rect 2668 13572 2724 13574
rect 2748 13572 2804 13574
rect 2828 13572 2884 13574
rect 2778 12724 2780 12744
rect 2780 12724 2832 12744
rect 2832 12724 2834 12744
rect 2778 12688 2834 12724
rect 2588 12538 2644 12540
rect 2668 12538 2724 12540
rect 2748 12538 2804 12540
rect 2828 12538 2884 12540
rect 2588 12486 2634 12538
rect 2634 12486 2644 12538
rect 2668 12486 2698 12538
rect 2698 12486 2710 12538
rect 2710 12486 2724 12538
rect 2748 12486 2762 12538
rect 2762 12486 2774 12538
rect 2774 12486 2804 12538
rect 2828 12486 2838 12538
rect 2838 12486 2884 12538
rect 2588 12484 2644 12486
rect 2668 12484 2724 12486
rect 2748 12484 2804 12486
rect 2828 12484 2884 12486
rect 2588 11450 2644 11452
rect 2668 11450 2724 11452
rect 2748 11450 2804 11452
rect 2828 11450 2884 11452
rect 2588 11398 2634 11450
rect 2634 11398 2644 11450
rect 2668 11398 2698 11450
rect 2698 11398 2710 11450
rect 2710 11398 2724 11450
rect 2748 11398 2762 11450
rect 2762 11398 2774 11450
rect 2774 11398 2804 11450
rect 2828 11398 2838 11450
rect 2838 11398 2884 11450
rect 2588 11396 2644 11398
rect 2668 11396 2724 11398
rect 2748 11396 2804 11398
rect 2828 11396 2884 11398
rect 2588 10362 2644 10364
rect 2668 10362 2724 10364
rect 2748 10362 2804 10364
rect 2828 10362 2884 10364
rect 2588 10310 2634 10362
rect 2634 10310 2644 10362
rect 2668 10310 2698 10362
rect 2698 10310 2710 10362
rect 2710 10310 2724 10362
rect 2748 10310 2762 10362
rect 2762 10310 2774 10362
rect 2774 10310 2804 10362
rect 2828 10310 2838 10362
rect 2838 10310 2884 10362
rect 2588 10308 2644 10310
rect 2668 10308 2724 10310
rect 2748 10308 2804 10310
rect 2828 10308 2884 10310
rect 2588 9274 2644 9276
rect 2668 9274 2724 9276
rect 2748 9274 2804 9276
rect 2828 9274 2884 9276
rect 2588 9222 2634 9274
rect 2634 9222 2644 9274
rect 2668 9222 2698 9274
rect 2698 9222 2710 9274
rect 2710 9222 2724 9274
rect 2748 9222 2762 9274
rect 2762 9222 2774 9274
rect 2774 9222 2804 9274
rect 2828 9222 2838 9274
rect 2838 9222 2884 9274
rect 2588 9220 2644 9222
rect 2668 9220 2724 9222
rect 2748 9220 2804 9222
rect 2828 9220 2884 9222
rect 2588 8186 2644 8188
rect 2668 8186 2724 8188
rect 2748 8186 2804 8188
rect 2828 8186 2884 8188
rect 2588 8134 2634 8186
rect 2634 8134 2644 8186
rect 2668 8134 2698 8186
rect 2698 8134 2710 8186
rect 2710 8134 2724 8186
rect 2748 8134 2762 8186
rect 2762 8134 2774 8186
rect 2774 8134 2804 8186
rect 2828 8134 2838 8186
rect 2838 8134 2884 8186
rect 2588 8132 2644 8134
rect 2668 8132 2724 8134
rect 2748 8132 2804 8134
rect 2828 8132 2884 8134
rect 2778 7248 2834 7304
rect 2588 7098 2644 7100
rect 2668 7098 2724 7100
rect 2748 7098 2804 7100
rect 2828 7098 2884 7100
rect 2588 7046 2634 7098
rect 2634 7046 2644 7098
rect 2668 7046 2698 7098
rect 2698 7046 2710 7098
rect 2710 7046 2724 7098
rect 2748 7046 2762 7098
rect 2762 7046 2774 7098
rect 2774 7046 2804 7098
rect 2828 7046 2838 7098
rect 2838 7046 2884 7098
rect 2588 7044 2644 7046
rect 2668 7044 2724 7046
rect 2748 7044 2804 7046
rect 2828 7044 2884 7046
rect 2588 6010 2644 6012
rect 2668 6010 2724 6012
rect 2748 6010 2804 6012
rect 2828 6010 2884 6012
rect 2588 5958 2634 6010
rect 2634 5958 2644 6010
rect 2668 5958 2698 6010
rect 2698 5958 2710 6010
rect 2710 5958 2724 6010
rect 2748 5958 2762 6010
rect 2762 5958 2774 6010
rect 2774 5958 2804 6010
rect 2828 5958 2838 6010
rect 2838 5958 2884 6010
rect 2588 5956 2644 5958
rect 2668 5956 2724 5958
rect 2748 5956 2804 5958
rect 2828 5956 2884 5958
rect 3238 15952 3294 16008
rect 3238 14864 3294 14920
rect 3422 19488 3478 19544
rect 4219 35930 4275 35932
rect 4299 35930 4355 35932
rect 4379 35930 4435 35932
rect 4459 35930 4515 35932
rect 4219 35878 4265 35930
rect 4265 35878 4275 35930
rect 4299 35878 4329 35930
rect 4329 35878 4341 35930
rect 4341 35878 4355 35930
rect 4379 35878 4393 35930
rect 4393 35878 4405 35930
rect 4405 35878 4435 35930
rect 4459 35878 4469 35930
rect 4469 35878 4515 35930
rect 4219 35876 4275 35878
rect 4299 35876 4355 35878
rect 4379 35876 4435 35878
rect 4459 35876 4515 35878
rect 4219 34842 4275 34844
rect 4299 34842 4355 34844
rect 4379 34842 4435 34844
rect 4459 34842 4515 34844
rect 4219 34790 4265 34842
rect 4265 34790 4275 34842
rect 4299 34790 4329 34842
rect 4329 34790 4341 34842
rect 4341 34790 4355 34842
rect 4379 34790 4393 34842
rect 4393 34790 4405 34842
rect 4405 34790 4435 34842
rect 4459 34790 4469 34842
rect 4469 34790 4515 34842
rect 4219 34788 4275 34790
rect 4299 34788 4355 34790
rect 4379 34788 4435 34790
rect 4459 34788 4515 34790
rect 4219 33754 4275 33756
rect 4299 33754 4355 33756
rect 4379 33754 4435 33756
rect 4459 33754 4515 33756
rect 4219 33702 4265 33754
rect 4265 33702 4275 33754
rect 4299 33702 4329 33754
rect 4329 33702 4341 33754
rect 4341 33702 4355 33754
rect 4379 33702 4393 33754
rect 4393 33702 4405 33754
rect 4405 33702 4435 33754
rect 4459 33702 4469 33754
rect 4469 33702 4515 33754
rect 4219 33700 4275 33702
rect 4299 33700 4355 33702
rect 4379 33700 4435 33702
rect 4459 33700 4515 33702
rect 4219 32666 4275 32668
rect 4299 32666 4355 32668
rect 4379 32666 4435 32668
rect 4459 32666 4515 32668
rect 4219 32614 4265 32666
rect 4265 32614 4275 32666
rect 4299 32614 4329 32666
rect 4329 32614 4341 32666
rect 4341 32614 4355 32666
rect 4379 32614 4393 32666
rect 4393 32614 4405 32666
rect 4405 32614 4435 32666
rect 4459 32614 4469 32666
rect 4469 32614 4515 32666
rect 4219 32612 4275 32614
rect 4299 32612 4355 32614
rect 4379 32612 4435 32614
rect 4459 32612 4515 32614
rect 4219 31578 4275 31580
rect 4299 31578 4355 31580
rect 4379 31578 4435 31580
rect 4459 31578 4515 31580
rect 4219 31526 4265 31578
rect 4265 31526 4275 31578
rect 4299 31526 4329 31578
rect 4329 31526 4341 31578
rect 4341 31526 4355 31578
rect 4379 31526 4393 31578
rect 4393 31526 4405 31578
rect 4405 31526 4435 31578
rect 4459 31526 4469 31578
rect 4469 31526 4515 31578
rect 4219 31524 4275 31526
rect 4299 31524 4355 31526
rect 4379 31524 4435 31526
rect 4459 31524 4515 31526
rect 4219 30490 4275 30492
rect 4299 30490 4355 30492
rect 4379 30490 4435 30492
rect 4459 30490 4515 30492
rect 4219 30438 4265 30490
rect 4265 30438 4275 30490
rect 4299 30438 4329 30490
rect 4329 30438 4341 30490
rect 4341 30438 4355 30490
rect 4379 30438 4393 30490
rect 4393 30438 4405 30490
rect 4405 30438 4435 30490
rect 4459 30438 4469 30490
rect 4469 30438 4515 30490
rect 4219 30436 4275 30438
rect 4299 30436 4355 30438
rect 4379 30436 4435 30438
rect 4459 30436 4515 30438
rect 4219 29402 4275 29404
rect 4299 29402 4355 29404
rect 4379 29402 4435 29404
rect 4459 29402 4515 29404
rect 4219 29350 4265 29402
rect 4265 29350 4275 29402
rect 4299 29350 4329 29402
rect 4329 29350 4341 29402
rect 4341 29350 4355 29402
rect 4379 29350 4393 29402
rect 4393 29350 4405 29402
rect 4405 29350 4435 29402
rect 4459 29350 4469 29402
rect 4469 29350 4515 29402
rect 4219 29348 4275 29350
rect 4299 29348 4355 29350
rect 4379 29348 4435 29350
rect 4459 29348 4515 29350
rect 4894 46144 4950 46200
rect 4802 41656 4858 41712
rect 4986 45056 5042 45112
rect 4894 39480 4950 39536
rect 5078 41928 5134 41984
rect 3974 27920 4030 27976
rect 3974 27512 4030 27568
rect 4219 28314 4275 28316
rect 4299 28314 4355 28316
rect 4379 28314 4435 28316
rect 4459 28314 4515 28316
rect 4219 28262 4265 28314
rect 4265 28262 4275 28314
rect 4299 28262 4329 28314
rect 4329 28262 4341 28314
rect 4341 28262 4355 28314
rect 4379 28262 4393 28314
rect 4393 28262 4405 28314
rect 4405 28262 4435 28314
rect 4459 28262 4469 28314
rect 4469 28262 4515 28314
rect 4219 28260 4275 28262
rect 4299 28260 4355 28262
rect 4379 28260 4435 28262
rect 4459 28260 4515 28262
rect 4219 27226 4275 27228
rect 4299 27226 4355 27228
rect 4379 27226 4435 27228
rect 4459 27226 4515 27228
rect 4219 27174 4265 27226
rect 4265 27174 4275 27226
rect 4299 27174 4329 27226
rect 4329 27174 4341 27226
rect 4341 27174 4355 27226
rect 4379 27174 4393 27226
rect 4393 27174 4405 27226
rect 4405 27174 4435 27226
rect 4459 27174 4469 27226
rect 4469 27174 4515 27226
rect 4219 27172 4275 27174
rect 4299 27172 4355 27174
rect 4379 27172 4435 27174
rect 4459 27172 4515 27174
rect 3606 15156 3662 15192
rect 3606 15136 3608 15156
rect 3608 15136 3660 15156
rect 3660 15136 3662 15156
rect 2588 4922 2644 4924
rect 2668 4922 2724 4924
rect 2748 4922 2804 4924
rect 2828 4922 2884 4924
rect 2588 4870 2634 4922
rect 2634 4870 2644 4922
rect 2668 4870 2698 4922
rect 2698 4870 2710 4922
rect 2710 4870 2724 4922
rect 2748 4870 2762 4922
rect 2762 4870 2774 4922
rect 2774 4870 2804 4922
rect 2828 4870 2838 4922
rect 2838 4870 2884 4922
rect 2588 4868 2644 4870
rect 2668 4868 2724 4870
rect 2748 4868 2804 4870
rect 2828 4868 2884 4870
rect 2962 4664 3018 4720
rect 3974 21664 4030 21720
rect 3882 20712 3938 20768
rect 4219 26138 4275 26140
rect 4299 26138 4355 26140
rect 4379 26138 4435 26140
rect 4459 26138 4515 26140
rect 4219 26086 4265 26138
rect 4265 26086 4275 26138
rect 4299 26086 4329 26138
rect 4329 26086 4341 26138
rect 4341 26086 4355 26138
rect 4379 26086 4393 26138
rect 4393 26086 4405 26138
rect 4405 26086 4435 26138
rect 4459 26086 4469 26138
rect 4469 26086 4515 26138
rect 4219 26084 4275 26086
rect 4299 26084 4355 26086
rect 4379 26084 4435 26086
rect 4459 26084 4515 26086
rect 4219 25050 4275 25052
rect 4299 25050 4355 25052
rect 4379 25050 4435 25052
rect 4459 25050 4515 25052
rect 4219 24998 4265 25050
rect 4265 24998 4275 25050
rect 4299 24998 4329 25050
rect 4329 24998 4341 25050
rect 4341 24998 4355 25050
rect 4379 24998 4393 25050
rect 4393 24998 4405 25050
rect 4405 24998 4435 25050
rect 4459 24998 4469 25050
rect 4469 24998 4515 25050
rect 4219 24996 4275 24998
rect 4299 24996 4355 24998
rect 4379 24996 4435 24998
rect 4459 24996 4515 24998
rect 4219 23962 4275 23964
rect 4299 23962 4355 23964
rect 4379 23962 4435 23964
rect 4459 23962 4515 23964
rect 4219 23910 4265 23962
rect 4265 23910 4275 23962
rect 4299 23910 4329 23962
rect 4329 23910 4341 23962
rect 4341 23910 4355 23962
rect 4379 23910 4393 23962
rect 4393 23910 4405 23962
rect 4405 23910 4435 23962
rect 4459 23910 4469 23962
rect 4469 23910 4515 23962
rect 4219 23908 4275 23910
rect 4299 23908 4355 23910
rect 4379 23908 4435 23910
rect 4459 23908 4515 23910
rect 4219 22874 4275 22876
rect 4299 22874 4355 22876
rect 4379 22874 4435 22876
rect 4459 22874 4515 22876
rect 4219 22822 4265 22874
rect 4265 22822 4275 22874
rect 4299 22822 4329 22874
rect 4329 22822 4341 22874
rect 4341 22822 4355 22874
rect 4379 22822 4393 22874
rect 4393 22822 4405 22874
rect 4405 22822 4435 22874
rect 4459 22822 4469 22874
rect 4469 22822 4515 22874
rect 4219 22820 4275 22822
rect 4299 22820 4355 22822
rect 4379 22820 4435 22822
rect 4459 22820 4515 22822
rect 4219 21786 4275 21788
rect 4299 21786 4355 21788
rect 4379 21786 4435 21788
rect 4459 21786 4515 21788
rect 4219 21734 4265 21786
rect 4265 21734 4275 21786
rect 4299 21734 4329 21786
rect 4329 21734 4341 21786
rect 4341 21734 4355 21786
rect 4379 21734 4393 21786
rect 4393 21734 4405 21786
rect 4405 21734 4435 21786
rect 4459 21734 4469 21786
rect 4469 21734 4515 21786
rect 4219 21732 4275 21734
rect 4299 21732 4355 21734
rect 4379 21732 4435 21734
rect 4459 21732 4515 21734
rect 4219 20698 4275 20700
rect 4299 20698 4355 20700
rect 4379 20698 4435 20700
rect 4459 20698 4515 20700
rect 4219 20646 4265 20698
rect 4265 20646 4275 20698
rect 4299 20646 4329 20698
rect 4329 20646 4341 20698
rect 4341 20646 4355 20698
rect 4379 20646 4393 20698
rect 4393 20646 4405 20698
rect 4405 20646 4435 20698
rect 4459 20646 4469 20698
rect 4469 20646 4515 20698
rect 4219 20644 4275 20646
rect 4299 20644 4355 20646
rect 4379 20644 4435 20646
rect 4459 20644 4515 20646
rect 3974 20304 4030 20360
rect 4066 19896 4122 19952
rect 4219 19610 4275 19612
rect 4299 19610 4355 19612
rect 4379 19610 4435 19612
rect 4459 19610 4515 19612
rect 4219 19558 4265 19610
rect 4265 19558 4275 19610
rect 4299 19558 4329 19610
rect 4329 19558 4341 19610
rect 4341 19558 4355 19610
rect 4379 19558 4393 19610
rect 4393 19558 4405 19610
rect 4405 19558 4435 19610
rect 4459 19558 4469 19610
rect 4469 19558 4515 19610
rect 4219 19556 4275 19558
rect 4299 19556 4355 19558
rect 4379 19556 4435 19558
rect 4459 19556 4515 19558
rect 4219 18522 4275 18524
rect 4299 18522 4355 18524
rect 4379 18522 4435 18524
rect 4459 18522 4515 18524
rect 4219 18470 4265 18522
rect 4265 18470 4275 18522
rect 4299 18470 4329 18522
rect 4329 18470 4341 18522
rect 4341 18470 4355 18522
rect 4379 18470 4393 18522
rect 4393 18470 4405 18522
rect 4405 18470 4435 18522
rect 4459 18470 4469 18522
rect 4469 18470 4515 18522
rect 4219 18468 4275 18470
rect 4299 18468 4355 18470
rect 4379 18468 4435 18470
rect 4459 18468 4515 18470
rect 4219 17434 4275 17436
rect 4299 17434 4355 17436
rect 4379 17434 4435 17436
rect 4459 17434 4515 17436
rect 4219 17382 4265 17434
rect 4265 17382 4275 17434
rect 4299 17382 4329 17434
rect 4329 17382 4341 17434
rect 4341 17382 4355 17434
rect 4379 17382 4393 17434
rect 4393 17382 4405 17434
rect 4405 17382 4435 17434
rect 4459 17382 4469 17434
rect 4469 17382 4515 17434
rect 4219 17380 4275 17382
rect 4299 17380 4355 17382
rect 4379 17380 4435 17382
rect 4459 17380 4515 17382
rect 4219 16346 4275 16348
rect 4299 16346 4355 16348
rect 4379 16346 4435 16348
rect 4459 16346 4515 16348
rect 4219 16294 4265 16346
rect 4265 16294 4275 16346
rect 4299 16294 4329 16346
rect 4329 16294 4341 16346
rect 4341 16294 4355 16346
rect 4379 16294 4393 16346
rect 4393 16294 4405 16346
rect 4405 16294 4435 16346
rect 4459 16294 4469 16346
rect 4469 16294 4515 16346
rect 4219 16292 4275 16294
rect 4299 16292 4355 16294
rect 4379 16292 4435 16294
rect 4459 16292 4515 16294
rect 3882 14864 3938 14920
rect 3974 13912 4030 13968
rect 4219 15258 4275 15260
rect 4299 15258 4355 15260
rect 4379 15258 4435 15260
rect 4459 15258 4515 15260
rect 4219 15206 4265 15258
rect 4265 15206 4275 15258
rect 4299 15206 4329 15258
rect 4329 15206 4341 15258
rect 4341 15206 4355 15258
rect 4379 15206 4393 15258
rect 4393 15206 4405 15258
rect 4405 15206 4435 15258
rect 4459 15206 4469 15258
rect 4469 15206 4515 15258
rect 4219 15204 4275 15206
rect 4299 15204 4355 15206
rect 4379 15204 4435 15206
rect 4459 15204 4515 15206
rect 4158 14356 4160 14376
rect 4160 14356 4212 14376
rect 4212 14356 4214 14376
rect 4158 14320 4214 14356
rect 4219 14170 4275 14172
rect 4299 14170 4355 14172
rect 4379 14170 4435 14172
rect 4459 14170 4515 14172
rect 4219 14118 4265 14170
rect 4265 14118 4275 14170
rect 4299 14118 4329 14170
rect 4329 14118 4341 14170
rect 4341 14118 4355 14170
rect 4379 14118 4393 14170
rect 4393 14118 4405 14170
rect 4405 14118 4435 14170
rect 4459 14118 4469 14170
rect 4469 14118 4515 14170
rect 4219 14116 4275 14118
rect 4299 14116 4355 14118
rect 4379 14116 4435 14118
rect 4459 14116 4515 14118
rect 4066 13368 4122 13424
rect 4219 13082 4275 13084
rect 4299 13082 4355 13084
rect 4379 13082 4435 13084
rect 4459 13082 4515 13084
rect 4219 13030 4265 13082
rect 4265 13030 4275 13082
rect 4299 13030 4329 13082
rect 4329 13030 4341 13082
rect 4341 13030 4355 13082
rect 4379 13030 4393 13082
rect 4393 13030 4405 13082
rect 4405 13030 4435 13082
rect 4459 13030 4469 13082
rect 4469 13030 4515 13082
rect 4219 13028 4275 13030
rect 4299 13028 4355 13030
rect 4379 13028 4435 13030
rect 4459 13028 4515 13030
rect 4219 11994 4275 11996
rect 4299 11994 4355 11996
rect 4379 11994 4435 11996
rect 4459 11994 4515 11996
rect 4219 11942 4265 11994
rect 4265 11942 4275 11994
rect 4299 11942 4329 11994
rect 4329 11942 4341 11994
rect 4341 11942 4355 11994
rect 4379 11942 4393 11994
rect 4393 11942 4405 11994
rect 4405 11942 4435 11994
rect 4459 11942 4469 11994
rect 4469 11942 4515 11994
rect 4219 11940 4275 11942
rect 4299 11940 4355 11942
rect 4379 11940 4435 11942
rect 4459 11940 4515 11942
rect 3790 8744 3846 8800
rect 4219 10906 4275 10908
rect 4299 10906 4355 10908
rect 4379 10906 4435 10908
rect 4459 10906 4515 10908
rect 4219 10854 4265 10906
rect 4265 10854 4275 10906
rect 4299 10854 4329 10906
rect 4329 10854 4341 10906
rect 4341 10854 4355 10906
rect 4379 10854 4393 10906
rect 4393 10854 4405 10906
rect 4405 10854 4435 10906
rect 4459 10854 4469 10906
rect 4469 10854 4515 10906
rect 4219 10852 4275 10854
rect 4299 10852 4355 10854
rect 4379 10852 4435 10854
rect 4459 10852 4515 10854
rect 4219 9818 4275 9820
rect 4299 9818 4355 9820
rect 4379 9818 4435 9820
rect 4459 9818 4515 9820
rect 4219 9766 4265 9818
rect 4265 9766 4275 9818
rect 4299 9766 4329 9818
rect 4329 9766 4341 9818
rect 4341 9766 4355 9818
rect 4379 9766 4393 9818
rect 4393 9766 4405 9818
rect 4405 9766 4435 9818
rect 4459 9766 4469 9818
rect 4469 9766 4515 9818
rect 4219 9764 4275 9766
rect 4299 9764 4355 9766
rect 4379 9764 4435 9766
rect 4459 9764 4515 9766
rect 4219 8730 4275 8732
rect 4299 8730 4355 8732
rect 4379 8730 4435 8732
rect 4459 8730 4515 8732
rect 4219 8678 4265 8730
rect 4265 8678 4275 8730
rect 4299 8678 4329 8730
rect 4329 8678 4341 8730
rect 4341 8678 4355 8730
rect 4379 8678 4393 8730
rect 4393 8678 4405 8730
rect 4405 8678 4435 8730
rect 4459 8678 4469 8730
rect 4469 8678 4515 8730
rect 4219 8676 4275 8678
rect 4299 8676 4355 8678
rect 4379 8676 4435 8678
rect 4459 8676 4515 8678
rect 3422 5752 3478 5808
rect 5170 39752 5226 39808
rect 5078 36352 5134 36408
rect 5851 73466 5907 73468
rect 5931 73466 5987 73468
rect 6011 73466 6067 73468
rect 6091 73466 6147 73468
rect 5851 73414 5897 73466
rect 5897 73414 5907 73466
rect 5931 73414 5961 73466
rect 5961 73414 5973 73466
rect 5973 73414 5987 73466
rect 6011 73414 6025 73466
rect 6025 73414 6037 73466
rect 6037 73414 6067 73466
rect 6091 73414 6101 73466
rect 6101 73414 6147 73466
rect 5851 73412 5907 73414
rect 5931 73412 5987 73414
rect 6011 73412 6067 73414
rect 6091 73412 6147 73414
rect 5851 72378 5907 72380
rect 5931 72378 5987 72380
rect 6011 72378 6067 72380
rect 6091 72378 6147 72380
rect 5851 72326 5897 72378
rect 5897 72326 5907 72378
rect 5931 72326 5961 72378
rect 5961 72326 5973 72378
rect 5973 72326 5987 72378
rect 6011 72326 6025 72378
rect 6025 72326 6037 72378
rect 6037 72326 6067 72378
rect 6091 72326 6101 72378
rect 6101 72326 6147 72378
rect 5851 72324 5907 72326
rect 5931 72324 5987 72326
rect 6011 72324 6067 72326
rect 6091 72324 6147 72326
rect 5851 71290 5907 71292
rect 5931 71290 5987 71292
rect 6011 71290 6067 71292
rect 6091 71290 6147 71292
rect 5851 71238 5897 71290
rect 5897 71238 5907 71290
rect 5931 71238 5961 71290
rect 5961 71238 5973 71290
rect 5973 71238 5987 71290
rect 6011 71238 6025 71290
rect 6025 71238 6037 71290
rect 6037 71238 6067 71290
rect 6091 71238 6101 71290
rect 6101 71238 6147 71290
rect 5851 71236 5907 71238
rect 5931 71236 5987 71238
rect 6011 71236 6067 71238
rect 6091 71236 6147 71238
rect 9115 75642 9171 75644
rect 9195 75642 9251 75644
rect 9275 75642 9331 75644
rect 9355 75642 9411 75644
rect 9115 75590 9161 75642
rect 9161 75590 9171 75642
rect 9195 75590 9225 75642
rect 9225 75590 9237 75642
rect 9237 75590 9251 75642
rect 9275 75590 9289 75642
rect 9289 75590 9301 75642
rect 9301 75590 9331 75642
rect 9355 75590 9365 75642
rect 9365 75590 9411 75642
rect 9115 75588 9171 75590
rect 9195 75588 9251 75590
rect 9275 75588 9331 75590
rect 9355 75588 9411 75590
rect 7483 75098 7539 75100
rect 7563 75098 7619 75100
rect 7643 75098 7699 75100
rect 7723 75098 7779 75100
rect 7483 75046 7529 75098
rect 7529 75046 7539 75098
rect 7563 75046 7593 75098
rect 7593 75046 7605 75098
rect 7605 75046 7619 75098
rect 7643 75046 7657 75098
rect 7657 75046 7669 75098
rect 7669 75046 7699 75098
rect 7723 75046 7733 75098
rect 7733 75046 7779 75098
rect 7483 75044 7539 75046
rect 7563 75044 7619 75046
rect 7643 75044 7699 75046
rect 7723 75044 7779 75046
rect 10138 76472 10194 76528
rect 10230 75656 10286 75712
rect 10138 74840 10194 74896
rect 7483 74010 7539 74012
rect 7563 74010 7619 74012
rect 7643 74010 7699 74012
rect 7723 74010 7779 74012
rect 7483 73958 7529 74010
rect 7529 73958 7539 74010
rect 7563 73958 7593 74010
rect 7593 73958 7605 74010
rect 7605 73958 7619 74010
rect 7643 73958 7657 74010
rect 7657 73958 7669 74010
rect 7669 73958 7699 74010
rect 7723 73958 7733 74010
rect 7733 73958 7779 74010
rect 7483 73956 7539 73958
rect 7563 73956 7619 73958
rect 7643 73956 7699 73958
rect 7723 73956 7779 73958
rect 7483 72922 7539 72924
rect 7563 72922 7619 72924
rect 7643 72922 7699 72924
rect 7723 72922 7779 72924
rect 7483 72870 7529 72922
rect 7529 72870 7539 72922
rect 7563 72870 7593 72922
rect 7593 72870 7605 72922
rect 7605 72870 7619 72922
rect 7643 72870 7657 72922
rect 7657 72870 7669 72922
rect 7669 72870 7699 72922
rect 7723 72870 7733 72922
rect 7733 72870 7779 72922
rect 7483 72868 7539 72870
rect 7563 72868 7619 72870
rect 7643 72868 7699 72870
rect 7723 72868 7779 72870
rect 7483 71834 7539 71836
rect 7563 71834 7619 71836
rect 7643 71834 7699 71836
rect 7723 71834 7779 71836
rect 7483 71782 7529 71834
rect 7529 71782 7539 71834
rect 7563 71782 7593 71834
rect 7593 71782 7605 71834
rect 7605 71782 7619 71834
rect 7643 71782 7657 71834
rect 7657 71782 7669 71834
rect 7669 71782 7699 71834
rect 7723 71782 7733 71834
rect 7733 71782 7779 71834
rect 7483 71780 7539 71782
rect 7563 71780 7619 71782
rect 7643 71780 7699 71782
rect 7723 71780 7779 71782
rect 7483 70746 7539 70748
rect 7563 70746 7619 70748
rect 7643 70746 7699 70748
rect 7723 70746 7779 70748
rect 7483 70694 7529 70746
rect 7529 70694 7539 70746
rect 7563 70694 7593 70746
rect 7593 70694 7605 70746
rect 7605 70694 7619 70746
rect 7643 70694 7657 70746
rect 7657 70694 7669 70746
rect 7669 70694 7699 70746
rect 7723 70694 7733 70746
rect 7733 70694 7779 70746
rect 7483 70692 7539 70694
rect 7563 70692 7619 70694
rect 7643 70692 7699 70694
rect 7723 70692 7779 70694
rect 5851 70202 5907 70204
rect 5931 70202 5987 70204
rect 6011 70202 6067 70204
rect 6091 70202 6147 70204
rect 5851 70150 5897 70202
rect 5897 70150 5907 70202
rect 5931 70150 5961 70202
rect 5961 70150 5973 70202
rect 5973 70150 5987 70202
rect 6011 70150 6025 70202
rect 6025 70150 6037 70202
rect 6037 70150 6067 70202
rect 6091 70150 6101 70202
rect 6101 70150 6147 70202
rect 5851 70148 5907 70150
rect 5931 70148 5987 70150
rect 6011 70148 6067 70150
rect 6091 70148 6147 70150
rect 5722 69436 5724 69456
rect 5724 69436 5776 69456
rect 5776 69436 5778 69456
rect 5722 69400 5778 69436
rect 5851 69114 5907 69116
rect 5931 69114 5987 69116
rect 6011 69114 6067 69116
rect 6091 69114 6147 69116
rect 5851 69062 5897 69114
rect 5897 69062 5907 69114
rect 5931 69062 5961 69114
rect 5961 69062 5973 69114
rect 5973 69062 5987 69114
rect 6011 69062 6025 69114
rect 6025 69062 6037 69114
rect 6037 69062 6067 69114
rect 6091 69062 6101 69114
rect 6101 69062 6147 69114
rect 5851 69060 5907 69062
rect 5931 69060 5987 69062
rect 6011 69060 6067 69062
rect 6091 69060 6147 69062
rect 5851 68026 5907 68028
rect 5931 68026 5987 68028
rect 6011 68026 6067 68028
rect 6091 68026 6147 68028
rect 5851 67974 5897 68026
rect 5897 67974 5907 68026
rect 5931 67974 5961 68026
rect 5961 67974 5973 68026
rect 5973 67974 5987 68026
rect 6011 67974 6025 68026
rect 6025 67974 6037 68026
rect 6037 67974 6067 68026
rect 6091 67974 6101 68026
rect 6101 67974 6147 68026
rect 5851 67972 5907 67974
rect 5931 67972 5987 67974
rect 6011 67972 6067 67974
rect 6091 67972 6147 67974
rect 5851 66938 5907 66940
rect 5931 66938 5987 66940
rect 6011 66938 6067 66940
rect 6091 66938 6147 66940
rect 5851 66886 5897 66938
rect 5897 66886 5907 66938
rect 5931 66886 5961 66938
rect 5961 66886 5973 66938
rect 5973 66886 5987 66938
rect 6011 66886 6025 66938
rect 6025 66886 6037 66938
rect 6037 66886 6067 66938
rect 6091 66886 6101 66938
rect 6101 66886 6147 66938
rect 5851 66884 5907 66886
rect 5931 66884 5987 66886
rect 6011 66884 6067 66886
rect 6091 66884 6147 66886
rect 5851 65850 5907 65852
rect 5931 65850 5987 65852
rect 6011 65850 6067 65852
rect 6091 65850 6147 65852
rect 5851 65798 5897 65850
rect 5897 65798 5907 65850
rect 5931 65798 5961 65850
rect 5961 65798 5973 65850
rect 5973 65798 5987 65850
rect 6011 65798 6025 65850
rect 6025 65798 6037 65850
rect 6037 65798 6067 65850
rect 6091 65798 6101 65850
rect 6101 65798 6147 65850
rect 5851 65796 5907 65798
rect 5931 65796 5987 65798
rect 6011 65796 6067 65798
rect 6091 65796 6147 65798
rect 5538 60696 5594 60752
rect 5851 64762 5907 64764
rect 5931 64762 5987 64764
rect 6011 64762 6067 64764
rect 6091 64762 6147 64764
rect 5851 64710 5897 64762
rect 5897 64710 5907 64762
rect 5931 64710 5961 64762
rect 5961 64710 5973 64762
rect 5973 64710 5987 64762
rect 6011 64710 6025 64762
rect 6025 64710 6037 64762
rect 6037 64710 6067 64762
rect 6091 64710 6101 64762
rect 6101 64710 6147 64762
rect 5851 64708 5907 64710
rect 5931 64708 5987 64710
rect 6011 64708 6067 64710
rect 6091 64708 6147 64710
rect 5851 63674 5907 63676
rect 5931 63674 5987 63676
rect 6011 63674 6067 63676
rect 6091 63674 6147 63676
rect 5851 63622 5897 63674
rect 5897 63622 5907 63674
rect 5931 63622 5961 63674
rect 5961 63622 5973 63674
rect 5973 63622 5987 63674
rect 6011 63622 6025 63674
rect 6025 63622 6037 63674
rect 6037 63622 6067 63674
rect 6091 63622 6101 63674
rect 6101 63622 6147 63674
rect 5851 63620 5907 63622
rect 5931 63620 5987 63622
rect 6011 63620 6067 63622
rect 6091 63620 6147 63622
rect 5851 62586 5907 62588
rect 5931 62586 5987 62588
rect 6011 62586 6067 62588
rect 6091 62586 6147 62588
rect 5851 62534 5897 62586
rect 5897 62534 5907 62586
rect 5931 62534 5961 62586
rect 5961 62534 5973 62586
rect 5973 62534 5987 62586
rect 6011 62534 6025 62586
rect 6025 62534 6037 62586
rect 6037 62534 6067 62586
rect 6091 62534 6101 62586
rect 6101 62534 6147 62586
rect 5851 62532 5907 62534
rect 5931 62532 5987 62534
rect 6011 62532 6067 62534
rect 6091 62532 6147 62534
rect 5851 61498 5907 61500
rect 5931 61498 5987 61500
rect 6011 61498 6067 61500
rect 6091 61498 6147 61500
rect 5851 61446 5897 61498
rect 5897 61446 5907 61498
rect 5931 61446 5961 61498
rect 5961 61446 5973 61498
rect 5973 61446 5987 61498
rect 6011 61446 6025 61498
rect 6025 61446 6037 61498
rect 6037 61446 6067 61498
rect 6091 61446 6101 61498
rect 6101 61446 6147 61498
rect 5851 61444 5907 61446
rect 5931 61444 5987 61446
rect 6011 61444 6067 61446
rect 6091 61444 6147 61446
rect 6182 60560 6238 60616
rect 5851 60410 5907 60412
rect 5931 60410 5987 60412
rect 6011 60410 6067 60412
rect 6091 60410 6147 60412
rect 5851 60358 5897 60410
rect 5897 60358 5907 60410
rect 5931 60358 5961 60410
rect 5961 60358 5973 60410
rect 5973 60358 5987 60410
rect 6011 60358 6025 60410
rect 6025 60358 6037 60410
rect 6037 60358 6067 60410
rect 6091 60358 6101 60410
rect 6101 60358 6147 60410
rect 5851 60356 5907 60358
rect 5931 60356 5987 60358
rect 6011 60356 6067 60358
rect 6091 60356 6147 60358
rect 5851 59322 5907 59324
rect 5931 59322 5987 59324
rect 6011 59322 6067 59324
rect 6091 59322 6147 59324
rect 5851 59270 5897 59322
rect 5897 59270 5907 59322
rect 5931 59270 5961 59322
rect 5961 59270 5973 59322
rect 5973 59270 5987 59322
rect 6011 59270 6025 59322
rect 6025 59270 6037 59322
rect 6037 59270 6067 59322
rect 6091 59270 6101 59322
rect 6101 59270 6147 59322
rect 5851 59268 5907 59270
rect 5931 59268 5987 59270
rect 6011 59268 6067 59270
rect 6091 59268 6147 59270
rect 5851 58234 5907 58236
rect 5931 58234 5987 58236
rect 6011 58234 6067 58236
rect 6091 58234 6147 58236
rect 5851 58182 5897 58234
rect 5897 58182 5907 58234
rect 5931 58182 5961 58234
rect 5961 58182 5973 58234
rect 5973 58182 5987 58234
rect 6011 58182 6025 58234
rect 6025 58182 6037 58234
rect 6037 58182 6067 58234
rect 6091 58182 6101 58234
rect 6101 58182 6147 58234
rect 5851 58180 5907 58182
rect 5931 58180 5987 58182
rect 6011 58180 6067 58182
rect 6091 58180 6147 58182
rect 5851 57146 5907 57148
rect 5931 57146 5987 57148
rect 6011 57146 6067 57148
rect 6091 57146 6147 57148
rect 5851 57094 5897 57146
rect 5897 57094 5907 57146
rect 5931 57094 5961 57146
rect 5961 57094 5973 57146
rect 5973 57094 5987 57146
rect 6011 57094 6025 57146
rect 6025 57094 6037 57146
rect 6037 57094 6067 57146
rect 6091 57094 6101 57146
rect 6101 57094 6147 57146
rect 5851 57092 5907 57094
rect 5931 57092 5987 57094
rect 6011 57092 6067 57094
rect 6091 57092 6147 57094
rect 5851 56058 5907 56060
rect 5931 56058 5987 56060
rect 6011 56058 6067 56060
rect 6091 56058 6147 56060
rect 5851 56006 5897 56058
rect 5897 56006 5907 56058
rect 5931 56006 5961 56058
rect 5961 56006 5973 56058
rect 5973 56006 5987 56058
rect 6011 56006 6025 56058
rect 6025 56006 6037 56058
rect 6037 56006 6067 56058
rect 6091 56006 6101 56058
rect 6101 56006 6147 56058
rect 5851 56004 5907 56006
rect 5931 56004 5987 56006
rect 6011 56004 6067 56006
rect 6091 56004 6147 56006
rect 5851 54970 5907 54972
rect 5931 54970 5987 54972
rect 6011 54970 6067 54972
rect 6091 54970 6147 54972
rect 5851 54918 5897 54970
rect 5897 54918 5907 54970
rect 5931 54918 5961 54970
rect 5961 54918 5973 54970
rect 5973 54918 5987 54970
rect 6011 54918 6025 54970
rect 6025 54918 6037 54970
rect 6037 54918 6067 54970
rect 6091 54918 6101 54970
rect 6101 54918 6147 54970
rect 5851 54916 5907 54918
rect 5931 54916 5987 54918
rect 6011 54916 6067 54918
rect 6091 54916 6147 54918
rect 5851 53882 5907 53884
rect 5931 53882 5987 53884
rect 6011 53882 6067 53884
rect 6091 53882 6147 53884
rect 5851 53830 5897 53882
rect 5897 53830 5907 53882
rect 5931 53830 5961 53882
rect 5961 53830 5973 53882
rect 5973 53830 5987 53882
rect 6011 53830 6025 53882
rect 6025 53830 6037 53882
rect 6037 53830 6067 53882
rect 6091 53830 6101 53882
rect 6101 53830 6147 53882
rect 5851 53828 5907 53830
rect 5931 53828 5987 53830
rect 6011 53828 6067 53830
rect 6091 53828 6147 53830
rect 5851 52794 5907 52796
rect 5931 52794 5987 52796
rect 6011 52794 6067 52796
rect 6091 52794 6147 52796
rect 5851 52742 5897 52794
rect 5897 52742 5907 52794
rect 5931 52742 5961 52794
rect 5961 52742 5973 52794
rect 5973 52742 5987 52794
rect 6011 52742 6025 52794
rect 6025 52742 6037 52794
rect 6037 52742 6067 52794
rect 6091 52742 6101 52794
rect 6101 52742 6147 52794
rect 5851 52740 5907 52742
rect 5931 52740 5987 52742
rect 6011 52740 6067 52742
rect 6091 52740 6147 52742
rect 5851 51706 5907 51708
rect 5931 51706 5987 51708
rect 6011 51706 6067 51708
rect 6091 51706 6147 51708
rect 5851 51654 5897 51706
rect 5897 51654 5907 51706
rect 5931 51654 5961 51706
rect 5961 51654 5973 51706
rect 5973 51654 5987 51706
rect 6011 51654 6025 51706
rect 6025 51654 6037 51706
rect 6037 51654 6067 51706
rect 6091 51654 6101 51706
rect 6101 51654 6147 51706
rect 5851 51652 5907 51654
rect 5931 51652 5987 51654
rect 6011 51652 6067 51654
rect 6091 51652 6147 51654
rect 5851 50618 5907 50620
rect 5931 50618 5987 50620
rect 6011 50618 6067 50620
rect 6091 50618 6147 50620
rect 5851 50566 5897 50618
rect 5897 50566 5907 50618
rect 5931 50566 5961 50618
rect 5961 50566 5973 50618
rect 5973 50566 5987 50618
rect 6011 50566 6025 50618
rect 6025 50566 6037 50618
rect 6037 50566 6067 50618
rect 6091 50566 6101 50618
rect 6101 50566 6147 50618
rect 5851 50564 5907 50566
rect 5931 50564 5987 50566
rect 6011 50564 6067 50566
rect 6091 50564 6147 50566
rect 5851 49530 5907 49532
rect 5931 49530 5987 49532
rect 6011 49530 6067 49532
rect 6091 49530 6147 49532
rect 5851 49478 5897 49530
rect 5897 49478 5907 49530
rect 5931 49478 5961 49530
rect 5961 49478 5973 49530
rect 5973 49478 5987 49530
rect 6011 49478 6025 49530
rect 6025 49478 6037 49530
rect 6037 49478 6067 49530
rect 6091 49478 6101 49530
rect 6101 49478 6147 49530
rect 5851 49476 5907 49478
rect 5931 49476 5987 49478
rect 6011 49476 6067 49478
rect 6091 49476 6147 49478
rect 5630 49000 5686 49056
rect 5538 48864 5594 48920
rect 5630 48456 5686 48512
rect 5538 48286 5594 48342
rect 5354 41520 5410 41576
rect 4986 35536 5042 35592
rect 5262 36352 5318 36408
rect 5851 48442 5907 48444
rect 5931 48442 5987 48444
rect 6011 48442 6067 48444
rect 6091 48442 6147 48444
rect 5851 48390 5897 48442
rect 5897 48390 5907 48442
rect 5931 48390 5961 48442
rect 5961 48390 5973 48442
rect 5973 48390 5987 48442
rect 6011 48390 6025 48442
rect 6025 48390 6037 48442
rect 6037 48390 6067 48442
rect 6091 48390 6101 48442
rect 6101 48390 6147 48442
rect 5851 48388 5907 48390
rect 5931 48388 5987 48390
rect 6011 48388 6067 48390
rect 6091 48388 6147 48390
rect 6182 47776 6238 47832
rect 5851 47354 5907 47356
rect 5931 47354 5987 47356
rect 6011 47354 6067 47356
rect 6091 47354 6147 47356
rect 5851 47302 5897 47354
rect 5897 47302 5907 47354
rect 5931 47302 5961 47354
rect 5961 47302 5973 47354
rect 5973 47302 5987 47354
rect 6011 47302 6025 47354
rect 6025 47302 6037 47354
rect 6037 47302 6067 47354
rect 6091 47302 6101 47354
rect 6101 47302 6147 47354
rect 5851 47300 5907 47302
rect 5931 47300 5987 47302
rect 6011 47300 6067 47302
rect 6091 47300 6147 47302
rect 5851 46266 5907 46268
rect 5931 46266 5987 46268
rect 6011 46266 6067 46268
rect 6091 46266 6147 46268
rect 5851 46214 5897 46266
rect 5897 46214 5907 46266
rect 5931 46214 5961 46266
rect 5961 46214 5973 46266
rect 5973 46214 5987 46266
rect 6011 46214 6025 46266
rect 6025 46214 6037 46266
rect 6037 46214 6067 46266
rect 6091 46214 6101 46266
rect 6101 46214 6147 46266
rect 5851 46212 5907 46214
rect 5931 46212 5987 46214
rect 6011 46212 6067 46214
rect 6091 46212 6147 46214
rect 5722 45872 5778 45928
rect 5851 45178 5907 45180
rect 5931 45178 5987 45180
rect 6011 45178 6067 45180
rect 6091 45178 6147 45180
rect 5851 45126 5897 45178
rect 5897 45126 5907 45178
rect 5931 45126 5961 45178
rect 5961 45126 5973 45178
rect 5973 45126 5987 45178
rect 6011 45126 6025 45178
rect 6025 45126 6037 45178
rect 6037 45126 6067 45178
rect 6091 45126 6101 45178
rect 6101 45126 6147 45178
rect 5851 45124 5907 45126
rect 5931 45124 5987 45126
rect 6011 45124 6067 45126
rect 6091 45124 6147 45126
rect 5851 44090 5907 44092
rect 5931 44090 5987 44092
rect 6011 44090 6067 44092
rect 6091 44090 6147 44092
rect 5851 44038 5897 44090
rect 5897 44038 5907 44090
rect 5931 44038 5961 44090
rect 5961 44038 5973 44090
rect 5973 44038 5987 44090
rect 6011 44038 6025 44090
rect 6025 44038 6037 44090
rect 6037 44038 6067 44090
rect 6091 44038 6101 44090
rect 6101 44038 6147 44090
rect 5851 44036 5907 44038
rect 5931 44036 5987 44038
rect 6011 44036 6067 44038
rect 6091 44036 6147 44038
rect 5851 43002 5907 43004
rect 5931 43002 5987 43004
rect 6011 43002 6067 43004
rect 6091 43002 6147 43004
rect 5851 42950 5897 43002
rect 5897 42950 5907 43002
rect 5931 42950 5961 43002
rect 5961 42950 5973 43002
rect 5973 42950 5987 43002
rect 6011 42950 6025 43002
rect 6025 42950 6037 43002
rect 6037 42950 6067 43002
rect 6091 42950 6101 43002
rect 6101 42950 6147 43002
rect 5851 42948 5907 42950
rect 5931 42948 5987 42950
rect 6011 42948 6067 42950
rect 6091 42948 6147 42950
rect 5851 41914 5907 41916
rect 5931 41914 5987 41916
rect 6011 41914 6067 41916
rect 6091 41914 6147 41916
rect 5851 41862 5897 41914
rect 5897 41862 5907 41914
rect 5931 41862 5961 41914
rect 5961 41862 5973 41914
rect 5973 41862 5987 41914
rect 6011 41862 6025 41914
rect 6025 41862 6037 41914
rect 6037 41862 6067 41914
rect 6091 41862 6101 41914
rect 6101 41862 6147 41914
rect 5851 41860 5907 41862
rect 5931 41860 5987 41862
rect 6011 41860 6067 41862
rect 6091 41860 6147 41862
rect 6182 41520 6238 41576
rect 5262 35128 5318 35184
rect 4219 7642 4275 7644
rect 4299 7642 4355 7644
rect 4379 7642 4435 7644
rect 4459 7642 4515 7644
rect 4219 7590 4265 7642
rect 4265 7590 4275 7642
rect 4299 7590 4329 7642
rect 4329 7590 4341 7642
rect 4341 7590 4355 7642
rect 4379 7590 4393 7642
rect 4393 7590 4405 7642
rect 4405 7590 4435 7642
rect 4459 7590 4469 7642
rect 4469 7590 4515 7642
rect 4219 7588 4275 7590
rect 4299 7588 4355 7590
rect 4379 7588 4435 7590
rect 4459 7588 4515 7590
rect 4219 6554 4275 6556
rect 4299 6554 4355 6556
rect 4379 6554 4435 6556
rect 4459 6554 4515 6556
rect 4219 6502 4265 6554
rect 4265 6502 4275 6554
rect 4299 6502 4329 6554
rect 4329 6502 4341 6554
rect 4341 6502 4355 6554
rect 4379 6502 4393 6554
rect 4393 6502 4405 6554
rect 4405 6502 4435 6554
rect 4459 6502 4469 6554
rect 4469 6502 4515 6554
rect 4219 6500 4275 6502
rect 4299 6500 4355 6502
rect 4379 6500 4435 6502
rect 4459 6500 4515 6502
rect 3790 6160 3846 6216
rect 2588 3834 2644 3836
rect 2668 3834 2724 3836
rect 2748 3834 2804 3836
rect 2828 3834 2884 3836
rect 2588 3782 2634 3834
rect 2634 3782 2644 3834
rect 2668 3782 2698 3834
rect 2698 3782 2710 3834
rect 2710 3782 2724 3834
rect 2748 3782 2762 3834
rect 2762 3782 2774 3834
rect 2774 3782 2804 3834
rect 2828 3782 2838 3834
rect 2838 3782 2884 3834
rect 2588 3780 2644 3782
rect 2668 3780 2724 3782
rect 2748 3780 2804 3782
rect 2828 3780 2884 3782
rect 2870 3576 2926 3632
rect 3606 3984 3662 4040
rect 2588 2746 2644 2748
rect 2668 2746 2724 2748
rect 2748 2746 2804 2748
rect 2828 2746 2884 2748
rect 2588 2694 2634 2746
rect 2634 2694 2644 2746
rect 2668 2694 2698 2746
rect 2698 2694 2710 2746
rect 2710 2694 2724 2746
rect 2748 2694 2762 2746
rect 2762 2694 2774 2746
rect 2774 2694 2804 2746
rect 2828 2694 2838 2746
rect 2838 2694 2884 2746
rect 2588 2692 2644 2694
rect 2668 2692 2724 2694
rect 2748 2692 2804 2694
rect 2828 2692 2884 2694
rect 3514 2216 3570 2272
rect 2870 1400 2926 1456
rect 4219 5466 4275 5468
rect 4299 5466 4355 5468
rect 4379 5466 4435 5468
rect 4459 5466 4515 5468
rect 4219 5414 4265 5466
rect 4265 5414 4275 5466
rect 4299 5414 4329 5466
rect 4329 5414 4341 5466
rect 4341 5414 4355 5466
rect 4379 5414 4393 5466
rect 4393 5414 4405 5466
rect 4405 5414 4435 5466
rect 4459 5414 4469 5466
rect 4469 5414 4515 5466
rect 4219 5412 4275 5414
rect 4299 5412 4355 5414
rect 4379 5412 4435 5414
rect 4459 5412 4515 5414
rect 3974 5208 4030 5264
rect 3974 4392 4030 4448
rect 4219 4378 4275 4380
rect 4299 4378 4355 4380
rect 4379 4378 4435 4380
rect 4459 4378 4515 4380
rect 4219 4326 4265 4378
rect 4265 4326 4275 4378
rect 4299 4326 4329 4378
rect 4329 4326 4341 4378
rect 4341 4326 4355 4378
rect 4379 4326 4393 4378
rect 4393 4326 4405 4378
rect 4405 4326 4435 4378
rect 4459 4326 4469 4378
rect 4469 4326 4515 4378
rect 4219 4324 4275 4326
rect 4299 4324 4355 4326
rect 4379 4324 4435 4326
rect 4459 4324 4515 4326
rect 5851 40826 5907 40828
rect 5931 40826 5987 40828
rect 6011 40826 6067 40828
rect 6091 40826 6147 40828
rect 5851 40774 5897 40826
rect 5897 40774 5907 40826
rect 5931 40774 5961 40826
rect 5961 40774 5973 40826
rect 5973 40774 5987 40826
rect 6011 40774 6025 40826
rect 6025 40774 6037 40826
rect 6037 40774 6067 40826
rect 6091 40774 6101 40826
rect 6101 40774 6147 40826
rect 5851 40772 5907 40774
rect 5931 40772 5987 40774
rect 6011 40772 6067 40774
rect 6091 40772 6147 40774
rect 5851 39738 5907 39740
rect 5931 39738 5987 39740
rect 6011 39738 6067 39740
rect 6091 39738 6147 39740
rect 5851 39686 5897 39738
rect 5897 39686 5907 39738
rect 5931 39686 5961 39738
rect 5961 39686 5973 39738
rect 5973 39686 5987 39738
rect 6011 39686 6025 39738
rect 6025 39686 6037 39738
rect 6037 39686 6067 39738
rect 6091 39686 6101 39738
rect 6101 39686 6147 39738
rect 5851 39684 5907 39686
rect 5931 39684 5987 39686
rect 6011 39684 6067 39686
rect 6091 39684 6147 39686
rect 5851 38650 5907 38652
rect 5931 38650 5987 38652
rect 6011 38650 6067 38652
rect 6091 38650 6147 38652
rect 5851 38598 5897 38650
rect 5897 38598 5907 38650
rect 5931 38598 5961 38650
rect 5961 38598 5973 38650
rect 5973 38598 5987 38650
rect 6011 38598 6025 38650
rect 6025 38598 6037 38650
rect 6037 38598 6067 38650
rect 6091 38598 6101 38650
rect 6101 38598 6147 38650
rect 5851 38596 5907 38598
rect 5931 38596 5987 38598
rect 6011 38596 6067 38598
rect 6091 38596 6147 38598
rect 5851 37562 5907 37564
rect 5931 37562 5987 37564
rect 6011 37562 6067 37564
rect 6091 37562 6147 37564
rect 5851 37510 5897 37562
rect 5897 37510 5907 37562
rect 5931 37510 5961 37562
rect 5961 37510 5973 37562
rect 5973 37510 5987 37562
rect 6011 37510 6025 37562
rect 6025 37510 6037 37562
rect 6037 37510 6067 37562
rect 6091 37510 6101 37562
rect 6101 37510 6147 37562
rect 5851 37508 5907 37510
rect 5931 37508 5987 37510
rect 6011 37508 6067 37510
rect 6091 37508 6147 37510
rect 5851 36474 5907 36476
rect 5931 36474 5987 36476
rect 6011 36474 6067 36476
rect 6091 36474 6147 36476
rect 5851 36422 5897 36474
rect 5897 36422 5907 36474
rect 5931 36422 5961 36474
rect 5961 36422 5973 36474
rect 5973 36422 5987 36474
rect 6011 36422 6025 36474
rect 6025 36422 6037 36474
rect 6037 36422 6067 36474
rect 6091 36422 6101 36474
rect 6101 36422 6147 36474
rect 5851 36420 5907 36422
rect 5931 36420 5987 36422
rect 6011 36420 6067 36422
rect 6091 36420 6147 36422
rect 5851 35386 5907 35388
rect 5931 35386 5987 35388
rect 6011 35386 6067 35388
rect 6091 35386 6147 35388
rect 5851 35334 5897 35386
rect 5897 35334 5907 35386
rect 5931 35334 5961 35386
rect 5961 35334 5973 35386
rect 5973 35334 5987 35386
rect 6011 35334 6025 35386
rect 6025 35334 6037 35386
rect 6037 35334 6067 35386
rect 6091 35334 6101 35386
rect 6101 35334 6147 35386
rect 5851 35332 5907 35334
rect 5931 35332 5987 35334
rect 6011 35332 6067 35334
rect 6091 35332 6147 35334
rect 5851 34298 5907 34300
rect 5931 34298 5987 34300
rect 6011 34298 6067 34300
rect 6091 34298 6147 34300
rect 5851 34246 5897 34298
rect 5897 34246 5907 34298
rect 5931 34246 5961 34298
rect 5961 34246 5973 34298
rect 5973 34246 5987 34298
rect 6011 34246 6025 34298
rect 6025 34246 6037 34298
rect 6037 34246 6067 34298
rect 6091 34246 6101 34298
rect 6101 34246 6147 34298
rect 5851 34244 5907 34246
rect 5931 34244 5987 34246
rect 6011 34244 6067 34246
rect 6091 34244 6147 34246
rect 5851 33210 5907 33212
rect 5931 33210 5987 33212
rect 6011 33210 6067 33212
rect 6091 33210 6147 33212
rect 5851 33158 5897 33210
rect 5897 33158 5907 33210
rect 5931 33158 5961 33210
rect 5961 33158 5973 33210
rect 5973 33158 5987 33210
rect 6011 33158 6025 33210
rect 6025 33158 6037 33210
rect 6037 33158 6067 33210
rect 6091 33158 6101 33210
rect 6101 33158 6147 33210
rect 5851 33156 5907 33158
rect 5931 33156 5987 33158
rect 6011 33156 6067 33158
rect 6091 33156 6147 33158
rect 5851 32122 5907 32124
rect 5931 32122 5987 32124
rect 6011 32122 6067 32124
rect 6091 32122 6147 32124
rect 5851 32070 5897 32122
rect 5897 32070 5907 32122
rect 5931 32070 5961 32122
rect 5961 32070 5973 32122
rect 5973 32070 5987 32122
rect 6011 32070 6025 32122
rect 6025 32070 6037 32122
rect 6037 32070 6067 32122
rect 6091 32070 6101 32122
rect 6101 32070 6147 32122
rect 5851 32068 5907 32070
rect 5931 32068 5987 32070
rect 6011 32068 6067 32070
rect 6091 32068 6147 32070
rect 5851 31034 5907 31036
rect 5931 31034 5987 31036
rect 6011 31034 6067 31036
rect 6091 31034 6147 31036
rect 5851 30982 5897 31034
rect 5897 30982 5907 31034
rect 5931 30982 5961 31034
rect 5961 30982 5973 31034
rect 5973 30982 5987 31034
rect 6011 30982 6025 31034
rect 6025 30982 6037 31034
rect 6037 30982 6067 31034
rect 6091 30982 6101 31034
rect 6101 30982 6147 31034
rect 5851 30980 5907 30982
rect 5931 30980 5987 30982
rect 6011 30980 6067 30982
rect 6091 30980 6147 30982
rect 5851 29946 5907 29948
rect 5931 29946 5987 29948
rect 6011 29946 6067 29948
rect 6091 29946 6147 29948
rect 5851 29894 5897 29946
rect 5897 29894 5907 29946
rect 5931 29894 5961 29946
rect 5961 29894 5973 29946
rect 5973 29894 5987 29946
rect 6011 29894 6025 29946
rect 6025 29894 6037 29946
rect 6037 29894 6067 29946
rect 6091 29894 6101 29946
rect 6101 29894 6147 29946
rect 5851 29892 5907 29894
rect 5931 29892 5987 29894
rect 6011 29892 6067 29894
rect 6091 29892 6147 29894
rect 5851 28858 5907 28860
rect 5931 28858 5987 28860
rect 6011 28858 6067 28860
rect 6091 28858 6147 28860
rect 5851 28806 5897 28858
rect 5897 28806 5907 28858
rect 5931 28806 5961 28858
rect 5961 28806 5973 28858
rect 5973 28806 5987 28858
rect 6011 28806 6025 28858
rect 6025 28806 6037 28858
rect 6037 28806 6067 28858
rect 6091 28806 6101 28858
rect 6101 28806 6147 28858
rect 5851 28804 5907 28806
rect 5931 28804 5987 28806
rect 6011 28804 6067 28806
rect 6091 28804 6147 28806
rect 5851 27770 5907 27772
rect 5931 27770 5987 27772
rect 6011 27770 6067 27772
rect 6091 27770 6147 27772
rect 5851 27718 5897 27770
rect 5897 27718 5907 27770
rect 5931 27718 5961 27770
rect 5961 27718 5973 27770
rect 5973 27718 5987 27770
rect 6011 27718 6025 27770
rect 6025 27718 6037 27770
rect 6037 27718 6067 27770
rect 6091 27718 6101 27770
rect 6101 27718 6147 27770
rect 5851 27716 5907 27718
rect 5931 27716 5987 27718
rect 6011 27716 6067 27718
rect 6091 27716 6147 27718
rect 5851 26682 5907 26684
rect 5931 26682 5987 26684
rect 6011 26682 6067 26684
rect 6091 26682 6147 26684
rect 5851 26630 5897 26682
rect 5897 26630 5907 26682
rect 5931 26630 5961 26682
rect 5961 26630 5973 26682
rect 5973 26630 5987 26682
rect 6011 26630 6025 26682
rect 6025 26630 6037 26682
rect 6037 26630 6067 26682
rect 6091 26630 6101 26682
rect 6101 26630 6147 26682
rect 5851 26628 5907 26630
rect 5931 26628 5987 26630
rect 6011 26628 6067 26630
rect 6091 26628 6147 26630
rect 5851 25594 5907 25596
rect 5931 25594 5987 25596
rect 6011 25594 6067 25596
rect 6091 25594 6147 25596
rect 5851 25542 5897 25594
rect 5897 25542 5907 25594
rect 5931 25542 5961 25594
rect 5961 25542 5973 25594
rect 5973 25542 5987 25594
rect 6011 25542 6025 25594
rect 6025 25542 6037 25594
rect 6037 25542 6067 25594
rect 6091 25542 6101 25594
rect 6101 25542 6147 25594
rect 5851 25540 5907 25542
rect 5931 25540 5987 25542
rect 6011 25540 6067 25542
rect 6091 25540 6147 25542
rect 5851 24506 5907 24508
rect 5931 24506 5987 24508
rect 6011 24506 6067 24508
rect 6091 24506 6147 24508
rect 5851 24454 5897 24506
rect 5897 24454 5907 24506
rect 5931 24454 5961 24506
rect 5961 24454 5973 24506
rect 5973 24454 5987 24506
rect 6011 24454 6025 24506
rect 6025 24454 6037 24506
rect 6037 24454 6067 24506
rect 6091 24454 6101 24506
rect 6101 24454 6147 24506
rect 5851 24452 5907 24454
rect 5931 24452 5987 24454
rect 6011 24452 6067 24454
rect 6091 24452 6147 24454
rect 5851 23418 5907 23420
rect 5931 23418 5987 23420
rect 6011 23418 6067 23420
rect 6091 23418 6147 23420
rect 5851 23366 5897 23418
rect 5897 23366 5907 23418
rect 5931 23366 5961 23418
rect 5961 23366 5973 23418
rect 5973 23366 5987 23418
rect 6011 23366 6025 23418
rect 6025 23366 6037 23418
rect 6037 23366 6067 23418
rect 6091 23366 6101 23418
rect 6101 23366 6147 23418
rect 5851 23364 5907 23366
rect 5931 23364 5987 23366
rect 6011 23364 6067 23366
rect 6091 23364 6147 23366
rect 5851 22330 5907 22332
rect 5931 22330 5987 22332
rect 6011 22330 6067 22332
rect 6091 22330 6147 22332
rect 5851 22278 5897 22330
rect 5897 22278 5907 22330
rect 5931 22278 5961 22330
rect 5961 22278 5973 22330
rect 5973 22278 5987 22330
rect 6011 22278 6025 22330
rect 6025 22278 6037 22330
rect 6037 22278 6067 22330
rect 6091 22278 6101 22330
rect 6101 22278 6147 22330
rect 5851 22276 5907 22278
rect 5931 22276 5987 22278
rect 6011 22276 6067 22278
rect 6091 22276 6147 22278
rect 5851 21242 5907 21244
rect 5931 21242 5987 21244
rect 6011 21242 6067 21244
rect 6091 21242 6147 21244
rect 5851 21190 5897 21242
rect 5897 21190 5907 21242
rect 5931 21190 5961 21242
rect 5961 21190 5973 21242
rect 5973 21190 5987 21242
rect 6011 21190 6025 21242
rect 6025 21190 6037 21242
rect 6037 21190 6067 21242
rect 6091 21190 6101 21242
rect 6101 21190 6147 21242
rect 5851 21188 5907 21190
rect 5931 21188 5987 21190
rect 6011 21188 6067 21190
rect 6091 21188 6147 21190
rect 5851 20154 5907 20156
rect 5931 20154 5987 20156
rect 6011 20154 6067 20156
rect 6091 20154 6147 20156
rect 5851 20102 5897 20154
rect 5897 20102 5907 20154
rect 5931 20102 5961 20154
rect 5961 20102 5973 20154
rect 5973 20102 5987 20154
rect 6011 20102 6025 20154
rect 6025 20102 6037 20154
rect 6037 20102 6067 20154
rect 6091 20102 6101 20154
rect 6101 20102 6147 20154
rect 5851 20100 5907 20102
rect 5931 20100 5987 20102
rect 6011 20100 6067 20102
rect 6091 20100 6147 20102
rect 5851 19066 5907 19068
rect 5931 19066 5987 19068
rect 6011 19066 6067 19068
rect 6091 19066 6147 19068
rect 5851 19014 5897 19066
rect 5897 19014 5907 19066
rect 5931 19014 5961 19066
rect 5961 19014 5973 19066
rect 5973 19014 5987 19066
rect 6011 19014 6025 19066
rect 6025 19014 6037 19066
rect 6037 19014 6067 19066
rect 6091 19014 6101 19066
rect 6101 19014 6147 19066
rect 5851 19012 5907 19014
rect 5931 19012 5987 19014
rect 6011 19012 6067 19014
rect 6091 19012 6147 19014
rect 5851 17978 5907 17980
rect 5931 17978 5987 17980
rect 6011 17978 6067 17980
rect 6091 17978 6147 17980
rect 5851 17926 5897 17978
rect 5897 17926 5907 17978
rect 5931 17926 5961 17978
rect 5961 17926 5973 17978
rect 5973 17926 5987 17978
rect 6011 17926 6025 17978
rect 6025 17926 6037 17978
rect 6037 17926 6067 17978
rect 6091 17926 6101 17978
rect 6101 17926 6147 17978
rect 5851 17924 5907 17926
rect 5931 17924 5987 17926
rect 6011 17924 6067 17926
rect 6091 17924 6147 17926
rect 5851 16890 5907 16892
rect 5931 16890 5987 16892
rect 6011 16890 6067 16892
rect 6091 16890 6147 16892
rect 5851 16838 5897 16890
rect 5897 16838 5907 16890
rect 5931 16838 5961 16890
rect 5961 16838 5973 16890
rect 5973 16838 5987 16890
rect 6011 16838 6025 16890
rect 6025 16838 6037 16890
rect 6037 16838 6067 16890
rect 6091 16838 6101 16890
rect 6101 16838 6147 16890
rect 5851 16836 5907 16838
rect 5931 16836 5987 16838
rect 6011 16836 6067 16838
rect 6091 16836 6147 16838
rect 5851 15802 5907 15804
rect 5931 15802 5987 15804
rect 6011 15802 6067 15804
rect 6091 15802 6147 15804
rect 5851 15750 5897 15802
rect 5897 15750 5907 15802
rect 5931 15750 5961 15802
rect 5961 15750 5973 15802
rect 5973 15750 5987 15802
rect 6011 15750 6025 15802
rect 6025 15750 6037 15802
rect 6037 15750 6067 15802
rect 6091 15750 6101 15802
rect 6101 15750 6147 15802
rect 5851 15748 5907 15750
rect 5931 15748 5987 15750
rect 6011 15748 6067 15750
rect 6091 15748 6147 15750
rect 5851 14714 5907 14716
rect 5931 14714 5987 14716
rect 6011 14714 6067 14716
rect 6091 14714 6147 14716
rect 5851 14662 5897 14714
rect 5897 14662 5907 14714
rect 5931 14662 5961 14714
rect 5961 14662 5973 14714
rect 5973 14662 5987 14714
rect 6011 14662 6025 14714
rect 6025 14662 6037 14714
rect 6037 14662 6067 14714
rect 6091 14662 6101 14714
rect 6101 14662 6147 14714
rect 5851 14660 5907 14662
rect 5931 14660 5987 14662
rect 6011 14660 6067 14662
rect 6091 14660 6147 14662
rect 5851 13626 5907 13628
rect 5931 13626 5987 13628
rect 6011 13626 6067 13628
rect 6091 13626 6147 13628
rect 5851 13574 5897 13626
rect 5897 13574 5907 13626
rect 5931 13574 5961 13626
rect 5961 13574 5973 13626
rect 5973 13574 5987 13626
rect 6011 13574 6025 13626
rect 6025 13574 6037 13626
rect 6037 13574 6067 13626
rect 6091 13574 6101 13626
rect 6101 13574 6147 13626
rect 5851 13572 5907 13574
rect 5931 13572 5987 13574
rect 6011 13572 6067 13574
rect 6091 13572 6147 13574
rect 5851 12538 5907 12540
rect 5931 12538 5987 12540
rect 6011 12538 6067 12540
rect 6091 12538 6147 12540
rect 5851 12486 5897 12538
rect 5897 12486 5907 12538
rect 5931 12486 5961 12538
rect 5961 12486 5973 12538
rect 5973 12486 5987 12538
rect 6011 12486 6025 12538
rect 6025 12486 6037 12538
rect 6037 12486 6067 12538
rect 6091 12486 6101 12538
rect 6101 12486 6147 12538
rect 5851 12484 5907 12486
rect 5931 12484 5987 12486
rect 6011 12484 6067 12486
rect 6091 12484 6147 12486
rect 6550 49136 6606 49192
rect 6458 46416 6514 46472
rect 6826 48592 6882 48648
rect 6274 27396 6330 27432
rect 6274 27376 6276 27396
rect 6276 27376 6328 27396
rect 6328 27376 6330 27396
rect 5851 11450 5907 11452
rect 5931 11450 5987 11452
rect 6011 11450 6067 11452
rect 6091 11450 6147 11452
rect 5851 11398 5897 11450
rect 5897 11398 5907 11450
rect 5931 11398 5961 11450
rect 5961 11398 5973 11450
rect 5973 11398 5987 11450
rect 6011 11398 6025 11450
rect 6025 11398 6037 11450
rect 6037 11398 6067 11450
rect 6091 11398 6101 11450
rect 6101 11398 6147 11450
rect 5851 11396 5907 11398
rect 5931 11396 5987 11398
rect 6011 11396 6067 11398
rect 6091 11396 6147 11398
rect 5851 10362 5907 10364
rect 5931 10362 5987 10364
rect 6011 10362 6067 10364
rect 6091 10362 6147 10364
rect 5851 10310 5897 10362
rect 5897 10310 5907 10362
rect 5931 10310 5961 10362
rect 5961 10310 5973 10362
rect 5973 10310 5987 10362
rect 6011 10310 6025 10362
rect 6025 10310 6037 10362
rect 6037 10310 6067 10362
rect 6091 10310 6101 10362
rect 6101 10310 6147 10362
rect 5851 10308 5907 10310
rect 5931 10308 5987 10310
rect 6011 10308 6067 10310
rect 6091 10308 6147 10310
rect 5851 9274 5907 9276
rect 5931 9274 5987 9276
rect 6011 9274 6067 9276
rect 6091 9274 6147 9276
rect 5851 9222 5897 9274
rect 5897 9222 5907 9274
rect 5931 9222 5961 9274
rect 5961 9222 5973 9274
rect 5973 9222 5987 9274
rect 6011 9222 6025 9274
rect 6025 9222 6037 9274
rect 6037 9222 6067 9274
rect 6091 9222 6101 9274
rect 6101 9222 6147 9274
rect 5851 9220 5907 9222
rect 5931 9220 5987 9222
rect 6011 9220 6067 9222
rect 6091 9220 6147 9222
rect 5851 8186 5907 8188
rect 5931 8186 5987 8188
rect 6011 8186 6067 8188
rect 6091 8186 6147 8188
rect 5851 8134 5897 8186
rect 5897 8134 5907 8186
rect 5931 8134 5961 8186
rect 5961 8134 5973 8186
rect 5973 8134 5987 8186
rect 6011 8134 6025 8186
rect 6025 8134 6037 8186
rect 6037 8134 6067 8186
rect 6091 8134 6101 8186
rect 6101 8134 6147 8186
rect 5851 8132 5907 8134
rect 5931 8132 5987 8134
rect 6011 8132 6067 8134
rect 6091 8132 6147 8134
rect 5851 7098 5907 7100
rect 5931 7098 5987 7100
rect 6011 7098 6067 7100
rect 6091 7098 6147 7100
rect 5851 7046 5897 7098
rect 5897 7046 5907 7098
rect 5931 7046 5961 7098
rect 5961 7046 5973 7098
rect 5973 7046 5987 7098
rect 6011 7046 6025 7098
rect 6025 7046 6037 7098
rect 6037 7046 6067 7098
rect 6091 7046 6101 7098
rect 6101 7046 6147 7098
rect 5851 7044 5907 7046
rect 5931 7044 5987 7046
rect 6011 7044 6067 7046
rect 6091 7044 6147 7046
rect 6458 41384 6514 41440
rect 5851 6010 5907 6012
rect 5931 6010 5987 6012
rect 6011 6010 6067 6012
rect 6091 6010 6147 6012
rect 5851 5958 5897 6010
rect 5897 5958 5907 6010
rect 5931 5958 5961 6010
rect 5961 5958 5973 6010
rect 5973 5958 5987 6010
rect 6011 5958 6025 6010
rect 6025 5958 6037 6010
rect 6037 5958 6067 6010
rect 6091 5958 6101 6010
rect 6101 5958 6147 6010
rect 5851 5956 5907 5958
rect 5931 5956 5987 5958
rect 6011 5956 6067 5958
rect 6091 5956 6147 5958
rect 5851 4922 5907 4924
rect 5931 4922 5987 4924
rect 6011 4922 6067 4924
rect 6091 4922 6147 4924
rect 5851 4870 5897 4922
rect 5897 4870 5907 4922
rect 5931 4870 5961 4922
rect 5961 4870 5973 4922
rect 5973 4870 5987 4922
rect 6011 4870 6025 4922
rect 6025 4870 6037 4922
rect 6037 4870 6067 4922
rect 6091 4870 6101 4922
rect 6101 4870 6147 4922
rect 5851 4868 5907 4870
rect 5931 4868 5987 4870
rect 6011 4868 6067 4870
rect 6091 4868 6147 4870
rect 6734 46008 6790 46064
rect 6734 41520 6790 41576
rect 6734 41248 6790 41304
rect 7483 69658 7539 69660
rect 7563 69658 7619 69660
rect 7643 69658 7699 69660
rect 7723 69658 7779 69660
rect 7483 69606 7529 69658
rect 7529 69606 7539 69658
rect 7563 69606 7593 69658
rect 7593 69606 7605 69658
rect 7605 69606 7619 69658
rect 7643 69606 7657 69658
rect 7657 69606 7669 69658
rect 7669 69606 7699 69658
rect 7723 69606 7733 69658
rect 7733 69606 7779 69658
rect 7483 69604 7539 69606
rect 7563 69604 7619 69606
rect 7643 69604 7699 69606
rect 7723 69604 7779 69606
rect 7483 68570 7539 68572
rect 7563 68570 7619 68572
rect 7643 68570 7699 68572
rect 7723 68570 7779 68572
rect 7483 68518 7529 68570
rect 7529 68518 7539 68570
rect 7563 68518 7593 68570
rect 7593 68518 7605 68570
rect 7605 68518 7619 68570
rect 7643 68518 7657 68570
rect 7657 68518 7669 68570
rect 7669 68518 7699 68570
rect 7723 68518 7733 68570
rect 7733 68518 7779 68570
rect 7483 68516 7539 68518
rect 7563 68516 7619 68518
rect 7643 68516 7699 68518
rect 7723 68516 7779 68518
rect 7010 46416 7066 46472
rect 7483 67482 7539 67484
rect 7563 67482 7619 67484
rect 7643 67482 7699 67484
rect 7723 67482 7779 67484
rect 7483 67430 7529 67482
rect 7529 67430 7539 67482
rect 7563 67430 7593 67482
rect 7593 67430 7605 67482
rect 7605 67430 7619 67482
rect 7643 67430 7657 67482
rect 7657 67430 7669 67482
rect 7669 67430 7699 67482
rect 7723 67430 7733 67482
rect 7733 67430 7779 67482
rect 7483 67428 7539 67430
rect 7563 67428 7619 67430
rect 7643 67428 7699 67430
rect 7723 67428 7779 67430
rect 7483 66394 7539 66396
rect 7563 66394 7619 66396
rect 7643 66394 7699 66396
rect 7723 66394 7779 66396
rect 7483 66342 7529 66394
rect 7529 66342 7539 66394
rect 7563 66342 7593 66394
rect 7593 66342 7605 66394
rect 7605 66342 7619 66394
rect 7643 66342 7657 66394
rect 7657 66342 7669 66394
rect 7669 66342 7699 66394
rect 7723 66342 7733 66394
rect 7733 66342 7779 66394
rect 7483 66340 7539 66342
rect 7563 66340 7619 66342
rect 7643 66340 7699 66342
rect 7723 66340 7779 66342
rect 7483 65306 7539 65308
rect 7563 65306 7619 65308
rect 7643 65306 7699 65308
rect 7723 65306 7779 65308
rect 7483 65254 7529 65306
rect 7529 65254 7539 65306
rect 7563 65254 7593 65306
rect 7593 65254 7605 65306
rect 7605 65254 7619 65306
rect 7643 65254 7657 65306
rect 7657 65254 7669 65306
rect 7669 65254 7699 65306
rect 7723 65254 7733 65306
rect 7733 65254 7779 65306
rect 7483 65252 7539 65254
rect 7563 65252 7619 65254
rect 7643 65252 7699 65254
rect 7723 65252 7779 65254
rect 7483 64218 7539 64220
rect 7563 64218 7619 64220
rect 7643 64218 7699 64220
rect 7723 64218 7779 64220
rect 7483 64166 7529 64218
rect 7529 64166 7539 64218
rect 7563 64166 7593 64218
rect 7593 64166 7605 64218
rect 7605 64166 7619 64218
rect 7643 64166 7657 64218
rect 7657 64166 7669 64218
rect 7669 64166 7699 64218
rect 7723 64166 7733 64218
rect 7733 64166 7779 64218
rect 7483 64164 7539 64166
rect 7563 64164 7619 64166
rect 7643 64164 7699 64166
rect 7723 64164 7779 64166
rect 7483 63130 7539 63132
rect 7563 63130 7619 63132
rect 7643 63130 7699 63132
rect 7723 63130 7779 63132
rect 7483 63078 7529 63130
rect 7529 63078 7539 63130
rect 7563 63078 7593 63130
rect 7593 63078 7605 63130
rect 7605 63078 7619 63130
rect 7643 63078 7657 63130
rect 7657 63078 7669 63130
rect 7669 63078 7699 63130
rect 7723 63078 7733 63130
rect 7733 63078 7779 63130
rect 7483 63076 7539 63078
rect 7563 63076 7619 63078
rect 7643 63076 7699 63078
rect 7723 63076 7779 63078
rect 7483 62042 7539 62044
rect 7563 62042 7619 62044
rect 7643 62042 7699 62044
rect 7723 62042 7779 62044
rect 7483 61990 7529 62042
rect 7529 61990 7539 62042
rect 7563 61990 7593 62042
rect 7593 61990 7605 62042
rect 7605 61990 7619 62042
rect 7643 61990 7657 62042
rect 7657 61990 7669 62042
rect 7669 61990 7699 62042
rect 7723 61990 7733 62042
rect 7733 61990 7779 62042
rect 7483 61988 7539 61990
rect 7563 61988 7619 61990
rect 7643 61988 7699 61990
rect 7723 61988 7779 61990
rect 7483 60954 7539 60956
rect 7563 60954 7619 60956
rect 7643 60954 7699 60956
rect 7723 60954 7779 60956
rect 7483 60902 7529 60954
rect 7529 60902 7539 60954
rect 7563 60902 7593 60954
rect 7593 60902 7605 60954
rect 7605 60902 7619 60954
rect 7643 60902 7657 60954
rect 7657 60902 7669 60954
rect 7669 60902 7699 60954
rect 7723 60902 7733 60954
rect 7733 60902 7779 60954
rect 7483 60900 7539 60902
rect 7563 60900 7619 60902
rect 7643 60900 7699 60902
rect 7723 60900 7779 60902
rect 7483 59866 7539 59868
rect 7563 59866 7619 59868
rect 7643 59866 7699 59868
rect 7723 59866 7779 59868
rect 7483 59814 7529 59866
rect 7529 59814 7539 59866
rect 7563 59814 7593 59866
rect 7593 59814 7605 59866
rect 7605 59814 7619 59866
rect 7643 59814 7657 59866
rect 7657 59814 7669 59866
rect 7669 59814 7699 59866
rect 7723 59814 7733 59866
rect 7733 59814 7779 59866
rect 7483 59812 7539 59814
rect 7563 59812 7619 59814
rect 7643 59812 7699 59814
rect 7723 59812 7779 59814
rect 7483 58778 7539 58780
rect 7563 58778 7619 58780
rect 7643 58778 7699 58780
rect 7723 58778 7779 58780
rect 7483 58726 7529 58778
rect 7529 58726 7539 58778
rect 7563 58726 7593 58778
rect 7593 58726 7605 58778
rect 7605 58726 7619 58778
rect 7643 58726 7657 58778
rect 7657 58726 7669 58778
rect 7669 58726 7699 58778
rect 7723 58726 7733 58778
rect 7733 58726 7779 58778
rect 7483 58724 7539 58726
rect 7563 58724 7619 58726
rect 7643 58724 7699 58726
rect 7723 58724 7779 58726
rect 7483 57690 7539 57692
rect 7563 57690 7619 57692
rect 7643 57690 7699 57692
rect 7723 57690 7779 57692
rect 7483 57638 7529 57690
rect 7529 57638 7539 57690
rect 7563 57638 7593 57690
rect 7593 57638 7605 57690
rect 7605 57638 7619 57690
rect 7643 57638 7657 57690
rect 7657 57638 7669 57690
rect 7669 57638 7699 57690
rect 7723 57638 7733 57690
rect 7733 57638 7779 57690
rect 7483 57636 7539 57638
rect 7563 57636 7619 57638
rect 7643 57636 7699 57638
rect 7723 57636 7779 57638
rect 7483 56602 7539 56604
rect 7563 56602 7619 56604
rect 7643 56602 7699 56604
rect 7723 56602 7779 56604
rect 7483 56550 7529 56602
rect 7529 56550 7539 56602
rect 7563 56550 7593 56602
rect 7593 56550 7605 56602
rect 7605 56550 7619 56602
rect 7643 56550 7657 56602
rect 7657 56550 7669 56602
rect 7669 56550 7699 56602
rect 7723 56550 7733 56602
rect 7733 56550 7779 56602
rect 7483 56548 7539 56550
rect 7563 56548 7619 56550
rect 7643 56548 7699 56550
rect 7723 56548 7779 56550
rect 7483 55514 7539 55516
rect 7563 55514 7619 55516
rect 7643 55514 7699 55516
rect 7723 55514 7779 55516
rect 7483 55462 7529 55514
rect 7529 55462 7539 55514
rect 7563 55462 7593 55514
rect 7593 55462 7605 55514
rect 7605 55462 7619 55514
rect 7643 55462 7657 55514
rect 7657 55462 7669 55514
rect 7669 55462 7699 55514
rect 7723 55462 7733 55514
rect 7733 55462 7779 55514
rect 7483 55460 7539 55462
rect 7563 55460 7619 55462
rect 7643 55460 7699 55462
rect 7723 55460 7779 55462
rect 7483 54426 7539 54428
rect 7563 54426 7619 54428
rect 7643 54426 7699 54428
rect 7723 54426 7779 54428
rect 7483 54374 7529 54426
rect 7529 54374 7539 54426
rect 7563 54374 7593 54426
rect 7593 54374 7605 54426
rect 7605 54374 7619 54426
rect 7643 54374 7657 54426
rect 7657 54374 7669 54426
rect 7669 54374 7699 54426
rect 7723 54374 7733 54426
rect 7733 54374 7779 54426
rect 7483 54372 7539 54374
rect 7563 54372 7619 54374
rect 7643 54372 7699 54374
rect 7723 54372 7779 54374
rect 7483 53338 7539 53340
rect 7563 53338 7619 53340
rect 7643 53338 7699 53340
rect 7723 53338 7779 53340
rect 7483 53286 7529 53338
rect 7529 53286 7539 53338
rect 7563 53286 7593 53338
rect 7593 53286 7605 53338
rect 7605 53286 7619 53338
rect 7643 53286 7657 53338
rect 7657 53286 7669 53338
rect 7669 53286 7699 53338
rect 7723 53286 7733 53338
rect 7733 53286 7779 53338
rect 7483 53284 7539 53286
rect 7563 53284 7619 53286
rect 7643 53284 7699 53286
rect 7723 53284 7779 53286
rect 7483 52250 7539 52252
rect 7563 52250 7619 52252
rect 7643 52250 7699 52252
rect 7723 52250 7779 52252
rect 7483 52198 7529 52250
rect 7529 52198 7539 52250
rect 7563 52198 7593 52250
rect 7593 52198 7605 52250
rect 7605 52198 7619 52250
rect 7643 52198 7657 52250
rect 7657 52198 7669 52250
rect 7669 52198 7699 52250
rect 7723 52198 7733 52250
rect 7733 52198 7779 52250
rect 7483 52196 7539 52198
rect 7563 52196 7619 52198
rect 7643 52196 7699 52198
rect 7723 52196 7779 52198
rect 7483 51162 7539 51164
rect 7563 51162 7619 51164
rect 7643 51162 7699 51164
rect 7723 51162 7779 51164
rect 7483 51110 7529 51162
rect 7529 51110 7539 51162
rect 7563 51110 7593 51162
rect 7593 51110 7605 51162
rect 7605 51110 7619 51162
rect 7643 51110 7657 51162
rect 7657 51110 7669 51162
rect 7669 51110 7699 51162
rect 7723 51110 7733 51162
rect 7733 51110 7779 51162
rect 7483 51108 7539 51110
rect 7563 51108 7619 51110
rect 7643 51108 7699 51110
rect 7723 51108 7779 51110
rect 7483 50074 7539 50076
rect 7563 50074 7619 50076
rect 7643 50074 7699 50076
rect 7723 50074 7779 50076
rect 7483 50022 7529 50074
rect 7529 50022 7539 50074
rect 7563 50022 7593 50074
rect 7593 50022 7605 50074
rect 7605 50022 7619 50074
rect 7643 50022 7657 50074
rect 7657 50022 7669 50074
rect 7669 50022 7699 50074
rect 7723 50022 7733 50074
rect 7733 50022 7779 50074
rect 7483 50020 7539 50022
rect 7563 50020 7619 50022
rect 7643 50020 7699 50022
rect 7723 50020 7779 50022
rect 7483 48986 7539 48988
rect 7563 48986 7619 48988
rect 7643 48986 7699 48988
rect 7723 48986 7779 48988
rect 7483 48934 7529 48986
rect 7529 48934 7539 48986
rect 7563 48934 7593 48986
rect 7593 48934 7605 48986
rect 7605 48934 7619 48986
rect 7643 48934 7657 48986
rect 7657 48934 7669 48986
rect 7669 48934 7699 48986
rect 7723 48934 7733 48986
rect 7733 48934 7779 48986
rect 7483 48932 7539 48934
rect 7563 48932 7619 48934
rect 7643 48932 7699 48934
rect 7723 48932 7779 48934
rect 7483 47898 7539 47900
rect 7563 47898 7619 47900
rect 7643 47898 7699 47900
rect 7723 47898 7779 47900
rect 7483 47846 7529 47898
rect 7529 47846 7539 47898
rect 7563 47846 7593 47898
rect 7593 47846 7605 47898
rect 7605 47846 7619 47898
rect 7643 47846 7657 47898
rect 7657 47846 7669 47898
rect 7669 47846 7699 47898
rect 7723 47846 7733 47898
rect 7733 47846 7779 47898
rect 7483 47844 7539 47846
rect 7563 47844 7619 47846
rect 7643 47844 7699 47846
rect 7723 47844 7779 47846
rect 7483 46810 7539 46812
rect 7563 46810 7619 46812
rect 7643 46810 7699 46812
rect 7723 46810 7779 46812
rect 7483 46758 7529 46810
rect 7529 46758 7539 46810
rect 7563 46758 7593 46810
rect 7593 46758 7605 46810
rect 7605 46758 7619 46810
rect 7643 46758 7657 46810
rect 7657 46758 7669 46810
rect 7669 46758 7699 46810
rect 7723 46758 7733 46810
rect 7733 46758 7779 46810
rect 7483 46756 7539 46758
rect 7563 46756 7619 46758
rect 7643 46756 7699 46758
rect 7723 46756 7779 46758
rect 7930 46416 7986 46472
rect 7483 45722 7539 45724
rect 7563 45722 7619 45724
rect 7643 45722 7699 45724
rect 7723 45722 7779 45724
rect 7483 45670 7529 45722
rect 7529 45670 7539 45722
rect 7563 45670 7593 45722
rect 7593 45670 7605 45722
rect 7605 45670 7619 45722
rect 7643 45670 7657 45722
rect 7657 45670 7669 45722
rect 7669 45670 7699 45722
rect 7723 45670 7733 45722
rect 7733 45670 7779 45722
rect 7483 45668 7539 45670
rect 7563 45668 7619 45670
rect 7643 45668 7699 45670
rect 7723 45668 7779 45670
rect 7483 44634 7539 44636
rect 7563 44634 7619 44636
rect 7643 44634 7699 44636
rect 7723 44634 7779 44636
rect 7483 44582 7529 44634
rect 7529 44582 7539 44634
rect 7563 44582 7593 44634
rect 7593 44582 7605 44634
rect 7605 44582 7619 44634
rect 7643 44582 7657 44634
rect 7657 44582 7669 44634
rect 7669 44582 7699 44634
rect 7723 44582 7733 44634
rect 7733 44582 7779 44634
rect 7483 44580 7539 44582
rect 7563 44580 7619 44582
rect 7643 44580 7699 44582
rect 7723 44580 7779 44582
rect 7483 43546 7539 43548
rect 7563 43546 7619 43548
rect 7643 43546 7699 43548
rect 7723 43546 7779 43548
rect 7483 43494 7529 43546
rect 7529 43494 7539 43546
rect 7563 43494 7593 43546
rect 7593 43494 7605 43546
rect 7605 43494 7619 43546
rect 7643 43494 7657 43546
rect 7657 43494 7669 43546
rect 7669 43494 7699 43546
rect 7723 43494 7733 43546
rect 7733 43494 7779 43546
rect 7483 43492 7539 43494
rect 7563 43492 7619 43494
rect 7643 43492 7699 43494
rect 7723 43492 7779 43494
rect 7483 42458 7539 42460
rect 7563 42458 7619 42460
rect 7643 42458 7699 42460
rect 7723 42458 7779 42460
rect 7483 42406 7529 42458
rect 7529 42406 7539 42458
rect 7563 42406 7593 42458
rect 7593 42406 7605 42458
rect 7605 42406 7619 42458
rect 7643 42406 7657 42458
rect 7657 42406 7669 42458
rect 7669 42406 7699 42458
rect 7723 42406 7733 42458
rect 7733 42406 7779 42458
rect 7483 42404 7539 42406
rect 7563 42404 7619 42406
rect 7643 42404 7699 42406
rect 7723 42404 7779 42406
rect 7483 41370 7539 41372
rect 7563 41370 7619 41372
rect 7643 41370 7699 41372
rect 7723 41370 7779 41372
rect 7483 41318 7529 41370
rect 7529 41318 7539 41370
rect 7563 41318 7593 41370
rect 7593 41318 7605 41370
rect 7605 41318 7619 41370
rect 7643 41318 7657 41370
rect 7657 41318 7669 41370
rect 7669 41318 7699 41370
rect 7723 41318 7733 41370
rect 7733 41318 7779 41370
rect 7483 41316 7539 41318
rect 7563 41316 7619 41318
rect 7643 41316 7699 41318
rect 7723 41316 7779 41318
rect 7483 40282 7539 40284
rect 7563 40282 7619 40284
rect 7643 40282 7699 40284
rect 7723 40282 7779 40284
rect 7483 40230 7529 40282
rect 7529 40230 7539 40282
rect 7563 40230 7593 40282
rect 7593 40230 7605 40282
rect 7605 40230 7619 40282
rect 7643 40230 7657 40282
rect 7657 40230 7669 40282
rect 7669 40230 7699 40282
rect 7723 40230 7733 40282
rect 7733 40230 7779 40282
rect 7483 40228 7539 40230
rect 7563 40228 7619 40230
rect 7643 40228 7699 40230
rect 7723 40228 7779 40230
rect 7483 39194 7539 39196
rect 7563 39194 7619 39196
rect 7643 39194 7699 39196
rect 7723 39194 7779 39196
rect 7483 39142 7529 39194
rect 7529 39142 7539 39194
rect 7563 39142 7593 39194
rect 7593 39142 7605 39194
rect 7605 39142 7619 39194
rect 7643 39142 7657 39194
rect 7657 39142 7669 39194
rect 7669 39142 7699 39194
rect 7723 39142 7733 39194
rect 7733 39142 7779 39194
rect 7483 39140 7539 39142
rect 7563 39140 7619 39142
rect 7643 39140 7699 39142
rect 7723 39140 7779 39142
rect 7483 38106 7539 38108
rect 7563 38106 7619 38108
rect 7643 38106 7699 38108
rect 7723 38106 7779 38108
rect 7483 38054 7529 38106
rect 7529 38054 7539 38106
rect 7563 38054 7593 38106
rect 7593 38054 7605 38106
rect 7605 38054 7619 38106
rect 7643 38054 7657 38106
rect 7657 38054 7669 38106
rect 7669 38054 7699 38106
rect 7723 38054 7733 38106
rect 7733 38054 7779 38106
rect 7483 38052 7539 38054
rect 7563 38052 7619 38054
rect 7643 38052 7699 38054
rect 7723 38052 7779 38054
rect 7483 37018 7539 37020
rect 7563 37018 7619 37020
rect 7643 37018 7699 37020
rect 7723 37018 7779 37020
rect 7483 36966 7529 37018
rect 7529 36966 7539 37018
rect 7563 36966 7593 37018
rect 7593 36966 7605 37018
rect 7605 36966 7619 37018
rect 7643 36966 7657 37018
rect 7657 36966 7669 37018
rect 7669 36966 7699 37018
rect 7723 36966 7733 37018
rect 7733 36966 7779 37018
rect 7483 36964 7539 36966
rect 7563 36964 7619 36966
rect 7643 36964 7699 36966
rect 7723 36964 7779 36966
rect 7483 35930 7539 35932
rect 7563 35930 7619 35932
rect 7643 35930 7699 35932
rect 7723 35930 7779 35932
rect 7483 35878 7529 35930
rect 7529 35878 7539 35930
rect 7563 35878 7593 35930
rect 7593 35878 7605 35930
rect 7605 35878 7619 35930
rect 7643 35878 7657 35930
rect 7657 35878 7669 35930
rect 7669 35878 7699 35930
rect 7723 35878 7733 35930
rect 7733 35878 7779 35930
rect 7483 35876 7539 35878
rect 7563 35876 7619 35878
rect 7643 35876 7699 35878
rect 7723 35876 7779 35878
rect 7483 34842 7539 34844
rect 7563 34842 7619 34844
rect 7643 34842 7699 34844
rect 7723 34842 7779 34844
rect 7483 34790 7529 34842
rect 7529 34790 7539 34842
rect 7563 34790 7593 34842
rect 7593 34790 7605 34842
rect 7605 34790 7619 34842
rect 7643 34790 7657 34842
rect 7657 34790 7669 34842
rect 7669 34790 7699 34842
rect 7723 34790 7733 34842
rect 7733 34790 7779 34842
rect 7483 34788 7539 34790
rect 7563 34788 7619 34790
rect 7643 34788 7699 34790
rect 7723 34788 7779 34790
rect 7483 33754 7539 33756
rect 7563 33754 7619 33756
rect 7643 33754 7699 33756
rect 7723 33754 7779 33756
rect 7483 33702 7529 33754
rect 7529 33702 7539 33754
rect 7563 33702 7593 33754
rect 7593 33702 7605 33754
rect 7605 33702 7619 33754
rect 7643 33702 7657 33754
rect 7657 33702 7669 33754
rect 7669 33702 7699 33754
rect 7723 33702 7733 33754
rect 7733 33702 7779 33754
rect 7483 33700 7539 33702
rect 7563 33700 7619 33702
rect 7643 33700 7699 33702
rect 7723 33700 7779 33702
rect 7483 32666 7539 32668
rect 7563 32666 7619 32668
rect 7643 32666 7699 32668
rect 7723 32666 7779 32668
rect 7483 32614 7529 32666
rect 7529 32614 7539 32666
rect 7563 32614 7593 32666
rect 7593 32614 7605 32666
rect 7605 32614 7619 32666
rect 7643 32614 7657 32666
rect 7657 32614 7669 32666
rect 7669 32614 7699 32666
rect 7723 32614 7733 32666
rect 7733 32614 7779 32666
rect 7483 32612 7539 32614
rect 7563 32612 7619 32614
rect 7643 32612 7699 32614
rect 7723 32612 7779 32614
rect 7483 31578 7539 31580
rect 7563 31578 7619 31580
rect 7643 31578 7699 31580
rect 7723 31578 7779 31580
rect 7483 31526 7529 31578
rect 7529 31526 7539 31578
rect 7563 31526 7593 31578
rect 7593 31526 7605 31578
rect 7605 31526 7619 31578
rect 7643 31526 7657 31578
rect 7657 31526 7669 31578
rect 7669 31526 7699 31578
rect 7723 31526 7733 31578
rect 7733 31526 7779 31578
rect 7483 31524 7539 31526
rect 7563 31524 7619 31526
rect 7643 31524 7699 31526
rect 7723 31524 7779 31526
rect 7483 30490 7539 30492
rect 7563 30490 7619 30492
rect 7643 30490 7699 30492
rect 7723 30490 7779 30492
rect 7483 30438 7529 30490
rect 7529 30438 7539 30490
rect 7563 30438 7593 30490
rect 7593 30438 7605 30490
rect 7605 30438 7619 30490
rect 7643 30438 7657 30490
rect 7657 30438 7669 30490
rect 7669 30438 7699 30490
rect 7723 30438 7733 30490
rect 7733 30438 7779 30490
rect 7483 30436 7539 30438
rect 7563 30436 7619 30438
rect 7643 30436 7699 30438
rect 7723 30436 7779 30438
rect 7483 29402 7539 29404
rect 7563 29402 7619 29404
rect 7643 29402 7699 29404
rect 7723 29402 7779 29404
rect 7483 29350 7529 29402
rect 7529 29350 7539 29402
rect 7563 29350 7593 29402
rect 7593 29350 7605 29402
rect 7605 29350 7619 29402
rect 7643 29350 7657 29402
rect 7657 29350 7669 29402
rect 7669 29350 7699 29402
rect 7723 29350 7733 29402
rect 7733 29350 7779 29402
rect 7483 29348 7539 29350
rect 7563 29348 7619 29350
rect 7643 29348 7699 29350
rect 7723 29348 7779 29350
rect 7483 28314 7539 28316
rect 7563 28314 7619 28316
rect 7643 28314 7699 28316
rect 7723 28314 7779 28316
rect 7483 28262 7529 28314
rect 7529 28262 7539 28314
rect 7563 28262 7593 28314
rect 7593 28262 7605 28314
rect 7605 28262 7619 28314
rect 7643 28262 7657 28314
rect 7657 28262 7669 28314
rect 7669 28262 7699 28314
rect 7723 28262 7733 28314
rect 7733 28262 7779 28314
rect 7483 28260 7539 28262
rect 7563 28260 7619 28262
rect 7643 28260 7699 28262
rect 7723 28260 7779 28262
rect 7483 27226 7539 27228
rect 7563 27226 7619 27228
rect 7643 27226 7699 27228
rect 7723 27226 7779 27228
rect 7483 27174 7529 27226
rect 7529 27174 7539 27226
rect 7563 27174 7593 27226
rect 7593 27174 7605 27226
rect 7605 27174 7619 27226
rect 7643 27174 7657 27226
rect 7657 27174 7669 27226
rect 7669 27174 7699 27226
rect 7723 27174 7733 27226
rect 7733 27174 7779 27226
rect 7483 27172 7539 27174
rect 7563 27172 7619 27174
rect 7643 27172 7699 27174
rect 7723 27172 7779 27174
rect 7483 26138 7539 26140
rect 7563 26138 7619 26140
rect 7643 26138 7699 26140
rect 7723 26138 7779 26140
rect 7483 26086 7529 26138
rect 7529 26086 7539 26138
rect 7563 26086 7593 26138
rect 7593 26086 7605 26138
rect 7605 26086 7619 26138
rect 7643 26086 7657 26138
rect 7657 26086 7669 26138
rect 7669 26086 7699 26138
rect 7723 26086 7733 26138
rect 7733 26086 7779 26138
rect 7483 26084 7539 26086
rect 7563 26084 7619 26086
rect 7643 26084 7699 26086
rect 7723 26084 7779 26086
rect 7483 25050 7539 25052
rect 7563 25050 7619 25052
rect 7643 25050 7699 25052
rect 7723 25050 7779 25052
rect 7483 24998 7529 25050
rect 7529 24998 7539 25050
rect 7563 24998 7593 25050
rect 7593 24998 7605 25050
rect 7605 24998 7619 25050
rect 7643 24998 7657 25050
rect 7657 24998 7669 25050
rect 7669 24998 7699 25050
rect 7723 24998 7733 25050
rect 7733 24998 7779 25050
rect 7483 24996 7539 24998
rect 7563 24996 7619 24998
rect 7643 24996 7699 24998
rect 7723 24996 7779 24998
rect 7483 23962 7539 23964
rect 7563 23962 7619 23964
rect 7643 23962 7699 23964
rect 7723 23962 7779 23964
rect 7483 23910 7529 23962
rect 7529 23910 7539 23962
rect 7563 23910 7593 23962
rect 7593 23910 7605 23962
rect 7605 23910 7619 23962
rect 7643 23910 7657 23962
rect 7657 23910 7669 23962
rect 7669 23910 7699 23962
rect 7723 23910 7733 23962
rect 7733 23910 7779 23962
rect 7483 23908 7539 23910
rect 7563 23908 7619 23910
rect 7643 23908 7699 23910
rect 7723 23908 7779 23910
rect 7483 22874 7539 22876
rect 7563 22874 7619 22876
rect 7643 22874 7699 22876
rect 7723 22874 7779 22876
rect 7483 22822 7529 22874
rect 7529 22822 7539 22874
rect 7563 22822 7593 22874
rect 7593 22822 7605 22874
rect 7605 22822 7619 22874
rect 7643 22822 7657 22874
rect 7657 22822 7669 22874
rect 7669 22822 7699 22874
rect 7723 22822 7733 22874
rect 7733 22822 7779 22874
rect 7483 22820 7539 22822
rect 7563 22820 7619 22822
rect 7643 22820 7699 22822
rect 7723 22820 7779 22822
rect 7483 21786 7539 21788
rect 7563 21786 7619 21788
rect 7643 21786 7699 21788
rect 7723 21786 7779 21788
rect 7483 21734 7529 21786
rect 7529 21734 7539 21786
rect 7563 21734 7593 21786
rect 7593 21734 7605 21786
rect 7605 21734 7619 21786
rect 7643 21734 7657 21786
rect 7657 21734 7669 21786
rect 7669 21734 7699 21786
rect 7723 21734 7733 21786
rect 7733 21734 7779 21786
rect 7483 21732 7539 21734
rect 7563 21732 7619 21734
rect 7643 21732 7699 21734
rect 7723 21732 7779 21734
rect 7483 20698 7539 20700
rect 7563 20698 7619 20700
rect 7643 20698 7699 20700
rect 7723 20698 7779 20700
rect 7483 20646 7529 20698
rect 7529 20646 7539 20698
rect 7563 20646 7593 20698
rect 7593 20646 7605 20698
rect 7605 20646 7619 20698
rect 7643 20646 7657 20698
rect 7657 20646 7669 20698
rect 7669 20646 7699 20698
rect 7723 20646 7733 20698
rect 7733 20646 7779 20698
rect 7483 20644 7539 20646
rect 7563 20644 7619 20646
rect 7643 20644 7699 20646
rect 7723 20644 7779 20646
rect 7483 19610 7539 19612
rect 7563 19610 7619 19612
rect 7643 19610 7699 19612
rect 7723 19610 7779 19612
rect 7483 19558 7529 19610
rect 7529 19558 7539 19610
rect 7563 19558 7593 19610
rect 7593 19558 7605 19610
rect 7605 19558 7619 19610
rect 7643 19558 7657 19610
rect 7657 19558 7669 19610
rect 7669 19558 7699 19610
rect 7723 19558 7733 19610
rect 7733 19558 7779 19610
rect 7483 19556 7539 19558
rect 7563 19556 7619 19558
rect 7643 19556 7699 19558
rect 7723 19556 7779 19558
rect 7483 18522 7539 18524
rect 7563 18522 7619 18524
rect 7643 18522 7699 18524
rect 7723 18522 7779 18524
rect 7483 18470 7529 18522
rect 7529 18470 7539 18522
rect 7563 18470 7593 18522
rect 7593 18470 7605 18522
rect 7605 18470 7619 18522
rect 7643 18470 7657 18522
rect 7657 18470 7669 18522
rect 7669 18470 7699 18522
rect 7723 18470 7733 18522
rect 7733 18470 7779 18522
rect 7483 18468 7539 18470
rect 7563 18468 7619 18470
rect 7643 18468 7699 18470
rect 7723 18468 7779 18470
rect 7483 17434 7539 17436
rect 7563 17434 7619 17436
rect 7643 17434 7699 17436
rect 7723 17434 7779 17436
rect 7483 17382 7529 17434
rect 7529 17382 7539 17434
rect 7563 17382 7593 17434
rect 7593 17382 7605 17434
rect 7605 17382 7619 17434
rect 7643 17382 7657 17434
rect 7657 17382 7669 17434
rect 7669 17382 7699 17434
rect 7723 17382 7733 17434
rect 7733 17382 7779 17434
rect 7483 17380 7539 17382
rect 7563 17380 7619 17382
rect 7643 17380 7699 17382
rect 7723 17380 7779 17382
rect 7483 16346 7539 16348
rect 7563 16346 7619 16348
rect 7643 16346 7699 16348
rect 7723 16346 7779 16348
rect 7483 16294 7529 16346
rect 7529 16294 7539 16346
rect 7563 16294 7593 16346
rect 7593 16294 7605 16346
rect 7605 16294 7619 16346
rect 7643 16294 7657 16346
rect 7657 16294 7669 16346
rect 7669 16294 7699 16346
rect 7723 16294 7733 16346
rect 7733 16294 7779 16346
rect 7483 16292 7539 16294
rect 7563 16292 7619 16294
rect 7643 16292 7699 16294
rect 7723 16292 7779 16294
rect 7483 15258 7539 15260
rect 7563 15258 7619 15260
rect 7643 15258 7699 15260
rect 7723 15258 7779 15260
rect 7483 15206 7529 15258
rect 7529 15206 7539 15258
rect 7563 15206 7593 15258
rect 7593 15206 7605 15258
rect 7605 15206 7619 15258
rect 7643 15206 7657 15258
rect 7657 15206 7669 15258
rect 7669 15206 7699 15258
rect 7723 15206 7733 15258
rect 7733 15206 7779 15258
rect 7483 15204 7539 15206
rect 7563 15204 7619 15206
rect 7643 15204 7699 15206
rect 7723 15204 7779 15206
rect 7483 14170 7539 14172
rect 7563 14170 7619 14172
rect 7643 14170 7699 14172
rect 7723 14170 7779 14172
rect 7483 14118 7529 14170
rect 7529 14118 7539 14170
rect 7563 14118 7593 14170
rect 7593 14118 7605 14170
rect 7605 14118 7619 14170
rect 7643 14118 7657 14170
rect 7657 14118 7669 14170
rect 7669 14118 7699 14170
rect 7723 14118 7733 14170
rect 7733 14118 7779 14170
rect 7483 14116 7539 14118
rect 7563 14116 7619 14118
rect 7643 14116 7699 14118
rect 7723 14116 7779 14118
rect 7483 13082 7539 13084
rect 7563 13082 7619 13084
rect 7643 13082 7699 13084
rect 7723 13082 7779 13084
rect 7483 13030 7529 13082
rect 7529 13030 7539 13082
rect 7563 13030 7593 13082
rect 7593 13030 7605 13082
rect 7605 13030 7619 13082
rect 7643 13030 7657 13082
rect 7657 13030 7669 13082
rect 7669 13030 7699 13082
rect 7723 13030 7733 13082
rect 7733 13030 7779 13082
rect 7483 13028 7539 13030
rect 7563 13028 7619 13030
rect 7643 13028 7699 13030
rect 7723 13028 7779 13030
rect 7930 36624 7986 36680
rect 8114 46008 8170 46064
rect 8114 36352 8170 36408
rect 7483 11994 7539 11996
rect 7563 11994 7619 11996
rect 7643 11994 7699 11996
rect 7723 11994 7779 11996
rect 7483 11942 7529 11994
rect 7529 11942 7539 11994
rect 7563 11942 7593 11994
rect 7593 11942 7605 11994
rect 7605 11942 7619 11994
rect 7643 11942 7657 11994
rect 7657 11942 7669 11994
rect 7669 11942 7699 11994
rect 7723 11942 7733 11994
rect 7733 11942 7779 11994
rect 7483 11940 7539 11942
rect 7563 11940 7619 11942
rect 7643 11940 7699 11942
rect 7723 11940 7779 11942
rect 7483 10906 7539 10908
rect 7563 10906 7619 10908
rect 7643 10906 7699 10908
rect 7723 10906 7779 10908
rect 7483 10854 7529 10906
rect 7529 10854 7539 10906
rect 7563 10854 7593 10906
rect 7593 10854 7605 10906
rect 7605 10854 7619 10906
rect 7643 10854 7657 10906
rect 7657 10854 7669 10906
rect 7669 10854 7699 10906
rect 7723 10854 7733 10906
rect 7733 10854 7779 10906
rect 7483 10852 7539 10854
rect 7563 10852 7619 10854
rect 7643 10852 7699 10854
rect 7723 10852 7779 10854
rect 7483 9818 7539 9820
rect 7563 9818 7619 9820
rect 7643 9818 7699 9820
rect 7723 9818 7779 9820
rect 7483 9766 7529 9818
rect 7529 9766 7539 9818
rect 7563 9766 7593 9818
rect 7593 9766 7605 9818
rect 7605 9766 7619 9818
rect 7643 9766 7657 9818
rect 7657 9766 7669 9818
rect 7669 9766 7699 9818
rect 7723 9766 7733 9818
rect 7733 9766 7779 9818
rect 7483 9764 7539 9766
rect 7563 9764 7619 9766
rect 7643 9764 7699 9766
rect 7723 9764 7779 9766
rect 7483 8730 7539 8732
rect 7563 8730 7619 8732
rect 7643 8730 7699 8732
rect 7723 8730 7779 8732
rect 7483 8678 7529 8730
rect 7529 8678 7539 8730
rect 7563 8678 7593 8730
rect 7593 8678 7605 8730
rect 7605 8678 7619 8730
rect 7643 8678 7657 8730
rect 7657 8678 7669 8730
rect 7669 8678 7699 8730
rect 7723 8678 7733 8730
rect 7733 8678 7779 8730
rect 7483 8676 7539 8678
rect 7563 8676 7619 8678
rect 7643 8676 7699 8678
rect 7723 8676 7779 8678
rect 7483 7642 7539 7644
rect 7563 7642 7619 7644
rect 7643 7642 7699 7644
rect 7723 7642 7779 7644
rect 7483 7590 7529 7642
rect 7529 7590 7539 7642
rect 7563 7590 7593 7642
rect 7593 7590 7605 7642
rect 7605 7590 7619 7642
rect 7643 7590 7657 7642
rect 7657 7590 7669 7642
rect 7669 7590 7699 7642
rect 7723 7590 7733 7642
rect 7733 7590 7779 7642
rect 7483 7588 7539 7590
rect 7563 7588 7619 7590
rect 7643 7588 7699 7590
rect 7723 7588 7779 7590
rect 7483 6554 7539 6556
rect 7563 6554 7619 6556
rect 7643 6554 7699 6556
rect 7723 6554 7779 6556
rect 7483 6502 7529 6554
rect 7529 6502 7539 6554
rect 7563 6502 7593 6554
rect 7593 6502 7605 6554
rect 7605 6502 7619 6554
rect 7643 6502 7657 6554
rect 7657 6502 7669 6554
rect 7669 6502 7699 6554
rect 7723 6502 7733 6554
rect 7733 6502 7779 6554
rect 7483 6500 7539 6502
rect 7563 6500 7619 6502
rect 7643 6500 7699 6502
rect 7723 6500 7779 6502
rect 7483 5466 7539 5468
rect 7563 5466 7619 5468
rect 7643 5466 7699 5468
rect 7723 5466 7779 5468
rect 7483 5414 7529 5466
rect 7529 5414 7539 5466
rect 7563 5414 7593 5466
rect 7593 5414 7605 5466
rect 7605 5414 7619 5466
rect 7643 5414 7657 5466
rect 7657 5414 7669 5466
rect 7669 5414 7699 5466
rect 7723 5414 7733 5466
rect 7733 5414 7779 5466
rect 7483 5412 7539 5414
rect 7563 5412 7619 5414
rect 7643 5412 7699 5414
rect 7723 5412 7779 5414
rect 5851 3834 5907 3836
rect 5931 3834 5987 3836
rect 6011 3834 6067 3836
rect 6091 3834 6147 3836
rect 5851 3782 5897 3834
rect 5897 3782 5907 3834
rect 5931 3782 5961 3834
rect 5961 3782 5973 3834
rect 5973 3782 5987 3834
rect 6011 3782 6025 3834
rect 6025 3782 6037 3834
rect 6037 3782 6067 3834
rect 6091 3782 6101 3834
rect 6101 3782 6147 3834
rect 5851 3780 5907 3782
rect 5931 3780 5987 3782
rect 6011 3780 6067 3782
rect 6091 3780 6147 3782
rect 4219 3290 4275 3292
rect 4299 3290 4355 3292
rect 4379 3290 4435 3292
rect 4459 3290 4515 3292
rect 4219 3238 4265 3290
rect 4265 3238 4275 3290
rect 4299 3238 4329 3290
rect 4329 3238 4341 3290
rect 4341 3238 4355 3290
rect 4379 3238 4393 3290
rect 4393 3238 4405 3290
rect 4405 3238 4435 3290
rect 4459 3238 4469 3290
rect 4469 3238 4515 3290
rect 4219 3236 4275 3238
rect 4299 3236 4355 3238
rect 4379 3236 4435 3238
rect 4459 3236 4515 3238
rect 7483 4378 7539 4380
rect 7563 4378 7619 4380
rect 7643 4378 7699 4380
rect 7723 4378 7779 4380
rect 7483 4326 7529 4378
rect 7529 4326 7539 4378
rect 7563 4326 7593 4378
rect 7593 4326 7605 4378
rect 7605 4326 7619 4378
rect 7643 4326 7657 4378
rect 7657 4326 7669 4378
rect 7669 4326 7699 4378
rect 7723 4326 7733 4378
rect 7733 4326 7779 4378
rect 7483 4324 7539 4326
rect 7563 4324 7619 4326
rect 7643 4324 7699 4326
rect 7723 4324 7779 4326
rect 9115 74554 9171 74556
rect 9195 74554 9251 74556
rect 9275 74554 9331 74556
rect 9355 74554 9411 74556
rect 9115 74502 9161 74554
rect 9161 74502 9171 74554
rect 9195 74502 9225 74554
rect 9225 74502 9237 74554
rect 9237 74502 9251 74554
rect 9275 74502 9289 74554
rect 9289 74502 9301 74554
rect 9301 74502 9331 74554
rect 9355 74502 9365 74554
rect 9365 74502 9411 74554
rect 9115 74500 9171 74502
rect 9195 74500 9251 74502
rect 9275 74500 9331 74502
rect 9355 74500 9411 74502
rect 10138 74196 10140 74216
rect 10140 74196 10192 74216
rect 10192 74196 10194 74216
rect 10138 74160 10194 74196
rect 9115 73466 9171 73468
rect 9195 73466 9251 73468
rect 9275 73466 9331 73468
rect 9355 73466 9411 73468
rect 9115 73414 9161 73466
rect 9161 73414 9171 73466
rect 9195 73414 9225 73466
rect 9225 73414 9237 73466
rect 9237 73414 9251 73466
rect 9275 73414 9289 73466
rect 9289 73414 9301 73466
rect 9301 73414 9331 73466
rect 9355 73414 9365 73466
rect 9365 73414 9411 73466
rect 9115 73412 9171 73414
rect 9195 73412 9251 73414
rect 9275 73412 9331 73414
rect 9355 73412 9411 73414
rect 9115 72378 9171 72380
rect 9195 72378 9251 72380
rect 9275 72378 9331 72380
rect 9355 72378 9411 72380
rect 9115 72326 9161 72378
rect 9161 72326 9171 72378
rect 9195 72326 9225 72378
rect 9225 72326 9237 72378
rect 9237 72326 9251 72378
rect 9275 72326 9289 72378
rect 9289 72326 9301 72378
rect 9301 72326 9331 72378
rect 9355 72326 9365 72378
rect 9365 72326 9411 72378
rect 9115 72324 9171 72326
rect 9195 72324 9251 72326
rect 9275 72324 9331 72326
rect 9355 72324 9411 72326
rect 10138 73344 10194 73400
rect 10138 72664 10194 72720
rect 9115 71290 9171 71292
rect 9195 71290 9251 71292
rect 9275 71290 9331 71292
rect 9355 71290 9411 71292
rect 9115 71238 9161 71290
rect 9161 71238 9171 71290
rect 9195 71238 9225 71290
rect 9225 71238 9237 71290
rect 9237 71238 9251 71290
rect 9275 71238 9289 71290
rect 9289 71238 9301 71290
rect 9301 71238 9331 71290
rect 9355 71238 9365 71290
rect 9365 71238 9411 71290
rect 9115 71236 9171 71238
rect 9195 71236 9251 71238
rect 9275 71236 9331 71238
rect 9355 71236 9411 71238
rect 10138 71848 10194 71904
rect 10138 71032 10194 71088
rect 10138 70352 10194 70408
rect 9115 70202 9171 70204
rect 9195 70202 9251 70204
rect 9275 70202 9331 70204
rect 9355 70202 9411 70204
rect 9115 70150 9161 70202
rect 9161 70150 9171 70202
rect 9195 70150 9225 70202
rect 9225 70150 9237 70202
rect 9237 70150 9251 70202
rect 9275 70150 9289 70202
rect 9289 70150 9301 70202
rect 9301 70150 9331 70202
rect 9355 70150 9365 70202
rect 9365 70150 9411 70202
rect 9115 70148 9171 70150
rect 9195 70148 9251 70150
rect 9275 70148 9331 70150
rect 9355 70148 9411 70150
rect 10138 69536 10194 69592
rect 9115 69114 9171 69116
rect 9195 69114 9251 69116
rect 9275 69114 9331 69116
rect 9355 69114 9411 69116
rect 9115 69062 9161 69114
rect 9161 69062 9171 69114
rect 9195 69062 9225 69114
rect 9225 69062 9237 69114
rect 9237 69062 9251 69114
rect 9275 69062 9289 69114
rect 9289 69062 9301 69114
rect 9301 69062 9331 69114
rect 9355 69062 9365 69114
rect 9365 69062 9411 69114
rect 9115 69060 9171 69062
rect 9195 69060 9251 69062
rect 9275 69060 9331 69062
rect 9355 69060 9411 69062
rect 10138 68856 10194 68912
rect 10138 68040 10194 68096
rect 9115 68026 9171 68028
rect 9195 68026 9251 68028
rect 9275 68026 9331 68028
rect 9355 68026 9411 68028
rect 9115 67974 9161 68026
rect 9161 67974 9171 68026
rect 9195 67974 9225 68026
rect 9225 67974 9237 68026
rect 9237 67974 9251 68026
rect 9275 67974 9289 68026
rect 9289 67974 9301 68026
rect 9301 67974 9331 68026
rect 9355 67974 9365 68026
rect 9365 67974 9411 68026
rect 9115 67972 9171 67974
rect 9195 67972 9251 67974
rect 9275 67972 9331 67974
rect 9355 67972 9411 67974
rect 10138 67224 10194 67280
rect 9115 66938 9171 66940
rect 9195 66938 9251 66940
rect 9275 66938 9331 66940
rect 9355 66938 9411 66940
rect 9115 66886 9161 66938
rect 9161 66886 9171 66938
rect 9195 66886 9225 66938
rect 9225 66886 9237 66938
rect 9237 66886 9251 66938
rect 9275 66886 9289 66938
rect 9289 66886 9301 66938
rect 9301 66886 9331 66938
rect 9355 66886 9365 66938
rect 9365 66886 9411 66938
rect 9115 66884 9171 66886
rect 9195 66884 9251 66886
rect 9275 66884 9331 66886
rect 9355 66884 9411 66886
rect 10138 66580 10140 66600
rect 10140 66580 10192 66600
rect 10192 66580 10194 66600
rect 10138 66544 10194 66580
rect 9115 65850 9171 65852
rect 9195 65850 9251 65852
rect 9275 65850 9331 65852
rect 9355 65850 9411 65852
rect 9115 65798 9161 65850
rect 9161 65798 9171 65850
rect 9195 65798 9225 65850
rect 9225 65798 9237 65850
rect 9237 65798 9251 65850
rect 9275 65798 9289 65850
rect 9289 65798 9301 65850
rect 9301 65798 9331 65850
rect 9355 65798 9365 65850
rect 9365 65798 9411 65850
rect 9115 65796 9171 65798
rect 9195 65796 9251 65798
rect 9275 65796 9331 65798
rect 9355 65796 9411 65798
rect 9115 64762 9171 64764
rect 9195 64762 9251 64764
rect 9275 64762 9331 64764
rect 9355 64762 9411 64764
rect 9115 64710 9161 64762
rect 9161 64710 9171 64762
rect 9195 64710 9225 64762
rect 9225 64710 9237 64762
rect 9237 64710 9251 64762
rect 9275 64710 9289 64762
rect 9289 64710 9301 64762
rect 9301 64710 9331 64762
rect 9355 64710 9365 64762
rect 9365 64710 9411 64762
rect 9115 64708 9171 64710
rect 9195 64708 9251 64710
rect 9275 64708 9331 64710
rect 9355 64708 9411 64710
rect 9115 63674 9171 63676
rect 9195 63674 9251 63676
rect 9275 63674 9331 63676
rect 9355 63674 9411 63676
rect 9115 63622 9161 63674
rect 9161 63622 9171 63674
rect 9195 63622 9225 63674
rect 9225 63622 9237 63674
rect 9237 63622 9251 63674
rect 9275 63622 9289 63674
rect 9289 63622 9301 63674
rect 9301 63622 9331 63674
rect 9355 63622 9365 63674
rect 9365 63622 9411 63674
rect 9115 63620 9171 63622
rect 9195 63620 9251 63622
rect 9275 63620 9331 63622
rect 9355 63620 9411 63622
rect 10138 65728 10194 65784
rect 10138 65048 10194 65104
rect 10138 64232 10194 64288
rect 10138 63416 10194 63472
rect 10138 62736 10194 62792
rect 9115 62586 9171 62588
rect 9195 62586 9251 62588
rect 9275 62586 9331 62588
rect 9355 62586 9411 62588
rect 9115 62534 9161 62586
rect 9161 62534 9171 62586
rect 9195 62534 9225 62586
rect 9225 62534 9237 62586
rect 9237 62534 9251 62586
rect 9275 62534 9289 62586
rect 9289 62534 9301 62586
rect 9301 62534 9331 62586
rect 9355 62534 9365 62586
rect 9365 62534 9411 62586
rect 9115 62532 9171 62534
rect 9195 62532 9251 62534
rect 9275 62532 9331 62534
rect 9355 62532 9411 62534
rect 9115 61498 9171 61500
rect 9195 61498 9251 61500
rect 9275 61498 9331 61500
rect 9355 61498 9411 61500
rect 9115 61446 9161 61498
rect 9161 61446 9171 61498
rect 9195 61446 9225 61498
rect 9225 61446 9237 61498
rect 9237 61446 9251 61498
rect 9275 61446 9289 61498
rect 9289 61446 9301 61498
rect 9301 61446 9331 61498
rect 9355 61446 9365 61498
rect 9365 61446 9411 61498
rect 9115 61444 9171 61446
rect 9195 61444 9251 61446
rect 9275 61444 9331 61446
rect 9355 61444 9411 61446
rect 9115 60410 9171 60412
rect 9195 60410 9251 60412
rect 9275 60410 9331 60412
rect 9355 60410 9411 60412
rect 9115 60358 9161 60410
rect 9161 60358 9171 60410
rect 9195 60358 9225 60410
rect 9225 60358 9237 60410
rect 9237 60358 9251 60410
rect 9275 60358 9289 60410
rect 9289 60358 9301 60410
rect 9301 60358 9331 60410
rect 9355 60358 9365 60410
rect 9365 60358 9411 60410
rect 9115 60356 9171 60358
rect 9195 60356 9251 60358
rect 9275 60356 9331 60358
rect 9355 60356 9411 60358
rect 10138 61920 10194 61976
rect 9115 59322 9171 59324
rect 9195 59322 9251 59324
rect 9275 59322 9331 59324
rect 9355 59322 9411 59324
rect 9115 59270 9161 59322
rect 9161 59270 9171 59322
rect 9195 59270 9225 59322
rect 9225 59270 9237 59322
rect 9237 59270 9251 59322
rect 9275 59270 9289 59322
rect 9289 59270 9301 59322
rect 9301 59270 9331 59322
rect 9355 59270 9365 59322
rect 9365 59270 9411 59322
rect 9115 59268 9171 59270
rect 9195 59268 9251 59270
rect 9275 59268 9331 59270
rect 9355 59268 9411 59270
rect 10138 61240 10194 61296
rect 10138 60424 10194 60480
rect 10138 59608 10194 59664
rect 10138 58964 10140 58984
rect 10140 58964 10192 58984
rect 10192 58964 10194 58984
rect 10138 58928 10194 58964
rect 9115 58234 9171 58236
rect 9195 58234 9251 58236
rect 9275 58234 9331 58236
rect 9355 58234 9411 58236
rect 9115 58182 9161 58234
rect 9161 58182 9171 58234
rect 9195 58182 9225 58234
rect 9225 58182 9237 58234
rect 9237 58182 9251 58234
rect 9275 58182 9289 58234
rect 9289 58182 9301 58234
rect 9301 58182 9331 58234
rect 9355 58182 9365 58234
rect 9365 58182 9411 58234
rect 9115 58180 9171 58182
rect 9195 58180 9251 58182
rect 9275 58180 9331 58182
rect 9355 58180 9411 58182
rect 10138 58112 10194 58168
rect 10138 57432 10194 57488
rect 9115 57146 9171 57148
rect 9195 57146 9251 57148
rect 9275 57146 9331 57148
rect 9355 57146 9411 57148
rect 9115 57094 9161 57146
rect 9161 57094 9171 57146
rect 9195 57094 9225 57146
rect 9225 57094 9237 57146
rect 9237 57094 9251 57146
rect 9275 57094 9289 57146
rect 9289 57094 9301 57146
rect 9301 57094 9331 57146
rect 9355 57094 9365 57146
rect 9365 57094 9411 57146
rect 9115 57092 9171 57094
rect 9195 57092 9251 57094
rect 9275 57092 9331 57094
rect 9355 57092 9411 57094
rect 10138 56616 10194 56672
rect 9115 56058 9171 56060
rect 9195 56058 9251 56060
rect 9275 56058 9331 56060
rect 9355 56058 9411 56060
rect 9115 56006 9161 56058
rect 9161 56006 9171 56058
rect 9195 56006 9225 56058
rect 9225 56006 9237 56058
rect 9237 56006 9251 56058
rect 9275 56006 9289 56058
rect 9289 56006 9301 56058
rect 9301 56006 9331 56058
rect 9355 56006 9365 56058
rect 9365 56006 9411 56058
rect 9115 56004 9171 56006
rect 9195 56004 9251 56006
rect 9275 56004 9331 56006
rect 9355 56004 9411 56006
rect 10138 55800 10194 55856
rect 10138 55120 10194 55176
rect 9115 54970 9171 54972
rect 9195 54970 9251 54972
rect 9275 54970 9331 54972
rect 9355 54970 9411 54972
rect 9115 54918 9161 54970
rect 9161 54918 9171 54970
rect 9195 54918 9225 54970
rect 9225 54918 9237 54970
rect 9237 54918 9251 54970
rect 9275 54918 9289 54970
rect 9289 54918 9301 54970
rect 9301 54918 9331 54970
rect 9355 54918 9365 54970
rect 9365 54918 9411 54970
rect 9115 54916 9171 54918
rect 9195 54916 9251 54918
rect 9275 54916 9331 54918
rect 9355 54916 9411 54918
rect 9115 53882 9171 53884
rect 9195 53882 9251 53884
rect 9275 53882 9331 53884
rect 9355 53882 9411 53884
rect 9115 53830 9161 53882
rect 9161 53830 9171 53882
rect 9195 53830 9225 53882
rect 9225 53830 9237 53882
rect 9237 53830 9251 53882
rect 9275 53830 9289 53882
rect 9289 53830 9301 53882
rect 9301 53830 9331 53882
rect 9355 53830 9365 53882
rect 9365 53830 9411 53882
rect 9115 53828 9171 53830
rect 9195 53828 9251 53830
rect 9275 53828 9331 53830
rect 9355 53828 9411 53830
rect 9115 52794 9171 52796
rect 9195 52794 9251 52796
rect 9275 52794 9331 52796
rect 9355 52794 9411 52796
rect 9115 52742 9161 52794
rect 9161 52742 9171 52794
rect 9195 52742 9225 52794
rect 9225 52742 9237 52794
rect 9237 52742 9251 52794
rect 9275 52742 9289 52794
rect 9289 52742 9301 52794
rect 9301 52742 9331 52794
rect 9355 52742 9365 52794
rect 9365 52742 9411 52794
rect 9115 52740 9171 52742
rect 9195 52740 9251 52742
rect 9275 52740 9331 52742
rect 9355 52740 9411 52742
rect 10138 54304 10194 54360
rect 10046 53624 10102 53680
rect 10046 52844 10048 52864
rect 10048 52844 10100 52864
rect 10100 52844 10102 52864
rect 10046 52808 10102 52844
rect 10046 51992 10102 52048
rect 9115 51706 9171 51708
rect 9195 51706 9251 51708
rect 9275 51706 9331 51708
rect 9355 51706 9411 51708
rect 9115 51654 9161 51706
rect 9161 51654 9171 51706
rect 9195 51654 9225 51706
rect 9225 51654 9237 51706
rect 9237 51654 9251 51706
rect 9275 51654 9289 51706
rect 9289 51654 9301 51706
rect 9301 51654 9331 51706
rect 9355 51654 9365 51706
rect 9365 51654 9411 51706
rect 9115 51652 9171 51654
rect 9195 51652 9251 51654
rect 9275 51652 9331 51654
rect 9355 51652 9411 51654
rect 9115 50618 9171 50620
rect 9195 50618 9251 50620
rect 9275 50618 9331 50620
rect 9355 50618 9411 50620
rect 9115 50566 9161 50618
rect 9161 50566 9171 50618
rect 9195 50566 9225 50618
rect 9225 50566 9237 50618
rect 9237 50566 9251 50618
rect 9275 50566 9289 50618
rect 9289 50566 9301 50618
rect 9301 50566 9331 50618
rect 9355 50566 9365 50618
rect 9365 50566 9411 50618
rect 9115 50564 9171 50566
rect 9195 50564 9251 50566
rect 9275 50564 9331 50566
rect 9355 50564 9411 50566
rect 10046 51312 10102 51368
rect 10046 50496 10102 50552
rect 10046 49816 10102 49872
rect 9115 49530 9171 49532
rect 9195 49530 9251 49532
rect 9275 49530 9331 49532
rect 9355 49530 9411 49532
rect 9115 49478 9161 49530
rect 9161 49478 9171 49530
rect 9195 49478 9225 49530
rect 9225 49478 9237 49530
rect 9237 49478 9251 49530
rect 9275 49478 9289 49530
rect 9289 49478 9301 49530
rect 9301 49478 9331 49530
rect 9355 49478 9365 49530
rect 9365 49478 9411 49530
rect 9115 49476 9171 49478
rect 9195 49476 9251 49478
rect 9275 49476 9331 49478
rect 9355 49476 9411 49478
rect 9115 48442 9171 48444
rect 9195 48442 9251 48444
rect 9275 48442 9331 48444
rect 9355 48442 9411 48444
rect 9115 48390 9161 48442
rect 9161 48390 9171 48442
rect 9195 48390 9225 48442
rect 9225 48390 9237 48442
rect 9237 48390 9251 48442
rect 9275 48390 9289 48442
rect 9289 48390 9301 48442
rect 9301 48390 9331 48442
rect 9355 48390 9365 48442
rect 9365 48390 9411 48442
rect 9115 48388 9171 48390
rect 9195 48388 9251 48390
rect 9275 48388 9331 48390
rect 9355 48388 9411 48390
rect 9115 47354 9171 47356
rect 9195 47354 9251 47356
rect 9275 47354 9331 47356
rect 9355 47354 9411 47356
rect 9115 47302 9161 47354
rect 9161 47302 9171 47354
rect 9195 47302 9225 47354
rect 9225 47302 9237 47354
rect 9237 47302 9251 47354
rect 9275 47302 9289 47354
rect 9289 47302 9301 47354
rect 9301 47302 9331 47354
rect 9355 47302 9365 47354
rect 9365 47302 9411 47354
rect 9115 47300 9171 47302
rect 9195 47300 9251 47302
rect 9275 47300 9331 47302
rect 9355 47300 9411 47302
rect 10046 49036 10048 49056
rect 10048 49036 10100 49056
rect 10100 49036 10102 49056
rect 10046 49000 10102 49036
rect 10046 48184 10102 48240
rect 10046 47524 10102 47560
rect 10046 47504 10048 47524
rect 10048 47504 10100 47524
rect 10100 47504 10102 47524
rect 10046 46688 10102 46744
rect 9115 46266 9171 46268
rect 9195 46266 9251 46268
rect 9275 46266 9331 46268
rect 9355 46266 9411 46268
rect 9115 46214 9161 46266
rect 9161 46214 9171 46266
rect 9195 46214 9225 46266
rect 9225 46214 9237 46266
rect 9237 46214 9251 46266
rect 9275 46214 9289 46266
rect 9289 46214 9301 46266
rect 9301 46214 9331 46266
rect 9355 46214 9365 46266
rect 9365 46214 9411 46266
rect 9115 46212 9171 46214
rect 9195 46212 9251 46214
rect 9275 46212 9331 46214
rect 9355 46212 9411 46214
rect 10046 46008 10102 46064
rect 10046 45228 10048 45248
rect 10048 45228 10100 45248
rect 10100 45228 10102 45248
rect 10046 45192 10102 45228
rect 9115 45178 9171 45180
rect 9195 45178 9251 45180
rect 9275 45178 9331 45180
rect 9355 45178 9411 45180
rect 9115 45126 9161 45178
rect 9161 45126 9171 45178
rect 9195 45126 9225 45178
rect 9225 45126 9237 45178
rect 9237 45126 9251 45178
rect 9275 45126 9289 45178
rect 9289 45126 9301 45178
rect 9301 45126 9331 45178
rect 9355 45126 9365 45178
rect 9365 45126 9411 45178
rect 9115 45124 9171 45126
rect 9195 45124 9251 45126
rect 9275 45124 9331 45126
rect 9355 45124 9411 45126
rect 9115 44090 9171 44092
rect 9195 44090 9251 44092
rect 9275 44090 9331 44092
rect 9355 44090 9411 44092
rect 9115 44038 9161 44090
rect 9161 44038 9171 44090
rect 9195 44038 9225 44090
rect 9225 44038 9237 44090
rect 9237 44038 9251 44090
rect 9275 44038 9289 44090
rect 9289 44038 9301 44090
rect 9301 44038 9331 44090
rect 9355 44038 9365 44090
rect 9365 44038 9411 44090
rect 9115 44036 9171 44038
rect 9195 44036 9251 44038
rect 9275 44036 9331 44038
rect 9355 44036 9411 44038
rect 10046 44376 10102 44432
rect 10046 43696 10102 43752
rect 9115 43002 9171 43004
rect 9195 43002 9251 43004
rect 9275 43002 9331 43004
rect 9355 43002 9411 43004
rect 9115 42950 9161 43002
rect 9161 42950 9171 43002
rect 9195 42950 9225 43002
rect 9225 42950 9237 43002
rect 9237 42950 9251 43002
rect 9275 42950 9289 43002
rect 9289 42950 9301 43002
rect 9301 42950 9331 43002
rect 9355 42950 9365 43002
rect 9365 42950 9411 43002
rect 9115 42948 9171 42950
rect 9195 42948 9251 42950
rect 9275 42948 9331 42950
rect 9355 42948 9411 42950
rect 10046 42880 10102 42936
rect 9115 41914 9171 41916
rect 9195 41914 9251 41916
rect 9275 41914 9331 41916
rect 9355 41914 9411 41916
rect 9115 41862 9161 41914
rect 9161 41862 9171 41914
rect 9195 41862 9225 41914
rect 9225 41862 9237 41914
rect 9237 41862 9251 41914
rect 9275 41862 9289 41914
rect 9289 41862 9301 41914
rect 9301 41862 9331 41914
rect 9355 41862 9365 41914
rect 9365 41862 9411 41914
rect 9115 41860 9171 41862
rect 9195 41860 9251 41862
rect 9275 41860 9331 41862
rect 9355 41860 9411 41862
rect 10046 42200 10102 42256
rect 10046 41420 10048 41440
rect 10048 41420 10100 41440
rect 10100 41420 10102 41440
rect 10046 41384 10102 41420
rect 9115 40826 9171 40828
rect 9195 40826 9251 40828
rect 9275 40826 9331 40828
rect 9355 40826 9411 40828
rect 9115 40774 9161 40826
rect 9161 40774 9171 40826
rect 9195 40774 9225 40826
rect 9225 40774 9237 40826
rect 9237 40774 9251 40826
rect 9275 40774 9289 40826
rect 9289 40774 9301 40826
rect 9301 40774 9331 40826
rect 9355 40774 9365 40826
rect 9365 40774 9411 40826
rect 9115 40772 9171 40774
rect 9195 40772 9251 40774
rect 9275 40772 9331 40774
rect 9355 40772 9411 40774
rect 9115 39738 9171 39740
rect 9195 39738 9251 39740
rect 9275 39738 9331 39740
rect 9355 39738 9411 39740
rect 9115 39686 9161 39738
rect 9161 39686 9171 39738
rect 9195 39686 9225 39738
rect 9225 39686 9237 39738
rect 9237 39686 9251 39738
rect 9275 39686 9289 39738
rect 9289 39686 9301 39738
rect 9301 39686 9331 39738
rect 9355 39686 9365 39738
rect 9365 39686 9411 39738
rect 9115 39684 9171 39686
rect 9195 39684 9251 39686
rect 9275 39684 9331 39686
rect 9355 39684 9411 39686
rect 10046 40568 10102 40624
rect 10046 39908 10102 39944
rect 10046 39888 10048 39908
rect 10048 39888 10100 39908
rect 10100 39888 10102 39908
rect 10046 39072 10102 39128
rect 9115 38650 9171 38652
rect 9195 38650 9251 38652
rect 9275 38650 9331 38652
rect 9355 38650 9411 38652
rect 9115 38598 9161 38650
rect 9161 38598 9171 38650
rect 9195 38598 9225 38650
rect 9225 38598 9237 38650
rect 9237 38598 9251 38650
rect 9275 38598 9289 38650
rect 9289 38598 9301 38650
rect 9301 38598 9331 38650
rect 9355 38598 9365 38650
rect 9365 38598 9411 38650
rect 9115 38596 9171 38598
rect 9195 38596 9251 38598
rect 9275 38596 9331 38598
rect 9355 38596 9411 38598
rect 10046 38392 10102 38448
rect 9115 37562 9171 37564
rect 9195 37562 9251 37564
rect 9275 37562 9331 37564
rect 9355 37562 9411 37564
rect 9115 37510 9161 37562
rect 9161 37510 9171 37562
rect 9195 37510 9225 37562
rect 9225 37510 9237 37562
rect 9237 37510 9251 37562
rect 9275 37510 9289 37562
rect 9289 37510 9301 37562
rect 9301 37510 9331 37562
rect 9355 37510 9365 37562
rect 9365 37510 9411 37562
rect 9115 37508 9171 37510
rect 9195 37508 9251 37510
rect 9275 37508 9331 37510
rect 9355 37508 9411 37510
rect 10046 37612 10048 37632
rect 10048 37612 10100 37632
rect 10100 37612 10102 37632
rect 10046 37576 10102 37612
rect 10046 36760 10102 36816
rect 9115 36474 9171 36476
rect 9195 36474 9251 36476
rect 9275 36474 9331 36476
rect 9355 36474 9411 36476
rect 9115 36422 9161 36474
rect 9161 36422 9171 36474
rect 9195 36422 9225 36474
rect 9225 36422 9237 36474
rect 9237 36422 9251 36474
rect 9275 36422 9289 36474
rect 9289 36422 9301 36474
rect 9301 36422 9331 36474
rect 9355 36422 9365 36474
rect 9365 36422 9411 36474
rect 9115 36420 9171 36422
rect 9195 36420 9251 36422
rect 9275 36420 9331 36422
rect 9355 36420 9411 36422
rect 9115 35386 9171 35388
rect 9195 35386 9251 35388
rect 9275 35386 9331 35388
rect 9355 35386 9411 35388
rect 9115 35334 9161 35386
rect 9161 35334 9171 35386
rect 9195 35334 9225 35386
rect 9225 35334 9237 35386
rect 9237 35334 9251 35386
rect 9275 35334 9289 35386
rect 9289 35334 9301 35386
rect 9301 35334 9331 35386
rect 9355 35334 9365 35386
rect 9365 35334 9411 35386
rect 9115 35332 9171 35334
rect 9195 35332 9251 35334
rect 9275 35332 9331 35334
rect 9355 35332 9411 35334
rect 9115 34298 9171 34300
rect 9195 34298 9251 34300
rect 9275 34298 9331 34300
rect 9355 34298 9411 34300
rect 9115 34246 9161 34298
rect 9161 34246 9171 34298
rect 9195 34246 9225 34298
rect 9225 34246 9237 34298
rect 9237 34246 9251 34298
rect 9275 34246 9289 34298
rect 9289 34246 9301 34298
rect 9301 34246 9331 34298
rect 9355 34246 9365 34298
rect 9365 34246 9411 34298
rect 9115 34244 9171 34246
rect 9195 34244 9251 34246
rect 9275 34244 9331 34246
rect 9355 34244 9411 34246
rect 9115 33210 9171 33212
rect 9195 33210 9251 33212
rect 9275 33210 9331 33212
rect 9355 33210 9411 33212
rect 9115 33158 9161 33210
rect 9161 33158 9171 33210
rect 9195 33158 9225 33210
rect 9225 33158 9237 33210
rect 9237 33158 9251 33210
rect 9275 33158 9289 33210
rect 9289 33158 9301 33210
rect 9301 33158 9331 33210
rect 9355 33158 9365 33210
rect 9365 33158 9411 33210
rect 9115 33156 9171 33158
rect 9195 33156 9251 33158
rect 9275 33156 9331 33158
rect 9355 33156 9411 33158
rect 10046 36080 10102 36136
rect 10046 35264 10102 35320
rect 10046 34584 10102 34640
rect 10046 33804 10048 33824
rect 10048 33804 10100 33824
rect 10100 33804 10102 33824
rect 10046 33768 10102 33804
rect 9115 32122 9171 32124
rect 9195 32122 9251 32124
rect 9275 32122 9331 32124
rect 9355 32122 9411 32124
rect 9115 32070 9161 32122
rect 9161 32070 9171 32122
rect 9195 32070 9225 32122
rect 9225 32070 9237 32122
rect 9237 32070 9251 32122
rect 9275 32070 9289 32122
rect 9289 32070 9301 32122
rect 9301 32070 9331 32122
rect 9355 32070 9365 32122
rect 9365 32070 9411 32122
rect 9115 32068 9171 32070
rect 9195 32068 9251 32070
rect 9275 32068 9331 32070
rect 9355 32068 9411 32070
rect 10046 32952 10102 33008
rect 10046 32292 10102 32328
rect 10046 32272 10048 32292
rect 10048 32272 10100 32292
rect 10100 32272 10102 32292
rect 10046 31456 10102 31512
rect 9115 31034 9171 31036
rect 9195 31034 9251 31036
rect 9275 31034 9331 31036
rect 9355 31034 9411 31036
rect 9115 30982 9161 31034
rect 9161 30982 9171 31034
rect 9195 30982 9225 31034
rect 9225 30982 9237 31034
rect 9237 30982 9251 31034
rect 9275 30982 9289 31034
rect 9289 30982 9301 31034
rect 9301 30982 9331 31034
rect 9355 30982 9365 31034
rect 9365 30982 9411 31034
rect 9115 30980 9171 30982
rect 9195 30980 9251 30982
rect 9275 30980 9331 30982
rect 9355 30980 9411 30982
rect 10046 30776 10102 30832
rect 9115 29946 9171 29948
rect 9195 29946 9251 29948
rect 9275 29946 9331 29948
rect 9355 29946 9411 29948
rect 9115 29894 9161 29946
rect 9161 29894 9171 29946
rect 9195 29894 9225 29946
rect 9225 29894 9237 29946
rect 9237 29894 9251 29946
rect 9275 29894 9289 29946
rect 9289 29894 9301 29946
rect 9301 29894 9331 29946
rect 9355 29894 9365 29946
rect 9365 29894 9411 29946
rect 9115 29892 9171 29894
rect 9195 29892 9251 29894
rect 9275 29892 9331 29894
rect 9355 29892 9411 29894
rect 9115 28858 9171 28860
rect 9195 28858 9251 28860
rect 9275 28858 9331 28860
rect 9355 28858 9411 28860
rect 9115 28806 9161 28858
rect 9161 28806 9171 28858
rect 9195 28806 9225 28858
rect 9225 28806 9237 28858
rect 9237 28806 9251 28858
rect 9275 28806 9289 28858
rect 9289 28806 9301 28858
rect 9301 28806 9331 28858
rect 9355 28806 9365 28858
rect 9365 28806 9411 28858
rect 9115 28804 9171 28806
rect 9195 28804 9251 28806
rect 9275 28804 9331 28806
rect 9355 28804 9411 28806
rect 9115 27770 9171 27772
rect 9195 27770 9251 27772
rect 9275 27770 9331 27772
rect 9355 27770 9411 27772
rect 9115 27718 9161 27770
rect 9161 27718 9171 27770
rect 9195 27718 9225 27770
rect 9225 27718 9237 27770
rect 9237 27718 9251 27770
rect 9275 27718 9289 27770
rect 9289 27718 9301 27770
rect 9301 27718 9331 27770
rect 9355 27718 9365 27770
rect 9365 27718 9411 27770
rect 9115 27716 9171 27718
rect 9195 27716 9251 27718
rect 9275 27716 9331 27718
rect 9355 27716 9411 27718
rect 10046 29996 10048 30016
rect 10048 29996 10100 30016
rect 10100 29996 10102 30016
rect 10046 29960 10102 29996
rect 10966 29180 10968 29200
rect 10968 29180 11020 29200
rect 11020 29180 11022 29200
rect 10966 29144 11022 29180
rect 10138 28464 10194 28520
rect 10138 27668 10194 27704
rect 10138 27648 10140 27668
rect 10140 27648 10192 27668
rect 10192 27648 10194 27668
rect 10138 26988 10194 27024
rect 10138 26968 10140 26988
rect 10140 26968 10192 26988
rect 10192 26968 10194 26988
rect 9115 26682 9171 26684
rect 9195 26682 9251 26684
rect 9275 26682 9331 26684
rect 9355 26682 9411 26684
rect 9115 26630 9161 26682
rect 9161 26630 9171 26682
rect 9195 26630 9225 26682
rect 9225 26630 9237 26682
rect 9237 26630 9251 26682
rect 9275 26630 9289 26682
rect 9289 26630 9301 26682
rect 9301 26630 9331 26682
rect 9355 26630 9365 26682
rect 9365 26630 9411 26682
rect 9115 26628 9171 26630
rect 9195 26628 9251 26630
rect 9275 26628 9331 26630
rect 9355 26628 9411 26630
rect 10138 26152 10194 26208
rect 9115 25594 9171 25596
rect 9195 25594 9251 25596
rect 9275 25594 9331 25596
rect 9355 25594 9411 25596
rect 9115 25542 9161 25594
rect 9161 25542 9171 25594
rect 9195 25542 9225 25594
rect 9225 25542 9237 25594
rect 9237 25542 9251 25594
rect 9275 25542 9289 25594
rect 9289 25542 9301 25594
rect 9301 25542 9331 25594
rect 9355 25542 9365 25594
rect 9365 25542 9411 25594
rect 9115 25540 9171 25542
rect 9195 25540 9251 25542
rect 9275 25540 9331 25542
rect 9355 25540 9411 25542
rect 10230 25336 10286 25392
rect 10138 24656 10194 24712
rect 9115 24506 9171 24508
rect 9195 24506 9251 24508
rect 9275 24506 9331 24508
rect 9355 24506 9411 24508
rect 9115 24454 9161 24506
rect 9161 24454 9171 24506
rect 9195 24454 9225 24506
rect 9225 24454 9237 24506
rect 9237 24454 9251 24506
rect 9275 24454 9289 24506
rect 9289 24454 9301 24506
rect 9301 24454 9331 24506
rect 9355 24454 9365 24506
rect 9365 24454 9411 24506
rect 9115 24452 9171 24454
rect 9195 24452 9251 24454
rect 9275 24452 9331 24454
rect 9355 24452 9411 24454
rect 10138 23840 10194 23896
rect 9115 23418 9171 23420
rect 9195 23418 9251 23420
rect 9275 23418 9331 23420
rect 9355 23418 9411 23420
rect 9115 23366 9161 23418
rect 9161 23366 9171 23418
rect 9195 23366 9225 23418
rect 9225 23366 9237 23418
rect 9237 23366 9251 23418
rect 9275 23366 9289 23418
rect 9289 23366 9301 23418
rect 9301 23366 9331 23418
rect 9355 23366 9365 23418
rect 9365 23366 9411 23418
rect 9115 23364 9171 23366
rect 9195 23364 9251 23366
rect 9275 23364 9331 23366
rect 9355 23364 9411 23366
rect 10046 23160 10102 23216
rect 9115 22330 9171 22332
rect 9195 22330 9251 22332
rect 9275 22330 9331 22332
rect 9355 22330 9411 22332
rect 9115 22278 9161 22330
rect 9161 22278 9171 22330
rect 9195 22278 9225 22330
rect 9225 22278 9237 22330
rect 9237 22278 9251 22330
rect 9275 22278 9289 22330
rect 9289 22278 9301 22330
rect 9301 22278 9331 22330
rect 9355 22278 9365 22330
rect 9365 22278 9411 22330
rect 9115 22276 9171 22278
rect 9195 22276 9251 22278
rect 9275 22276 9331 22278
rect 9355 22276 9411 22278
rect 9115 21242 9171 21244
rect 9195 21242 9251 21244
rect 9275 21242 9331 21244
rect 9355 21242 9411 21244
rect 9115 21190 9161 21242
rect 9161 21190 9171 21242
rect 9195 21190 9225 21242
rect 9225 21190 9237 21242
rect 9237 21190 9251 21242
rect 9275 21190 9289 21242
rect 9289 21190 9301 21242
rect 9301 21190 9331 21242
rect 9355 21190 9365 21242
rect 9365 21190 9411 21242
rect 9115 21188 9171 21190
rect 9195 21188 9251 21190
rect 9275 21188 9331 21190
rect 9355 21188 9411 21190
rect 9115 20154 9171 20156
rect 9195 20154 9251 20156
rect 9275 20154 9331 20156
rect 9355 20154 9411 20156
rect 9115 20102 9161 20154
rect 9161 20102 9171 20154
rect 9195 20102 9225 20154
rect 9225 20102 9237 20154
rect 9237 20102 9251 20154
rect 9275 20102 9289 20154
rect 9289 20102 9301 20154
rect 9301 20102 9331 20154
rect 9355 20102 9365 20154
rect 9365 20102 9411 20154
rect 9115 20100 9171 20102
rect 9195 20100 9251 20102
rect 9275 20100 9331 20102
rect 9355 20100 9411 20102
rect 9115 19066 9171 19068
rect 9195 19066 9251 19068
rect 9275 19066 9331 19068
rect 9355 19066 9411 19068
rect 9115 19014 9161 19066
rect 9161 19014 9171 19066
rect 9195 19014 9225 19066
rect 9225 19014 9237 19066
rect 9237 19014 9251 19066
rect 9275 19014 9289 19066
rect 9289 19014 9301 19066
rect 9301 19014 9331 19066
rect 9355 19014 9365 19066
rect 9365 19014 9411 19066
rect 9115 19012 9171 19014
rect 9195 19012 9251 19014
rect 9275 19012 9331 19014
rect 9355 19012 9411 19014
rect 10046 22380 10048 22400
rect 10048 22380 10100 22400
rect 10100 22380 10102 22400
rect 10046 22344 10102 22380
rect 9115 17978 9171 17980
rect 9195 17978 9251 17980
rect 9275 17978 9331 17980
rect 9355 17978 9411 17980
rect 9115 17926 9161 17978
rect 9161 17926 9171 17978
rect 9195 17926 9225 17978
rect 9225 17926 9237 17978
rect 9237 17926 9251 17978
rect 9275 17926 9289 17978
rect 9289 17926 9301 17978
rect 9301 17926 9331 17978
rect 9355 17926 9365 17978
rect 9365 17926 9411 17978
rect 9115 17924 9171 17926
rect 9195 17924 9251 17926
rect 9275 17924 9331 17926
rect 9355 17924 9411 17926
rect 9115 16890 9171 16892
rect 9195 16890 9251 16892
rect 9275 16890 9331 16892
rect 9355 16890 9411 16892
rect 9115 16838 9161 16890
rect 9161 16838 9171 16890
rect 9195 16838 9225 16890
rect 9225 16838 9237 16890
rect 9237 16838 9251 16890
rect 9275 16838 9289 16890
rect 9289 16838 9301 16890
rect 9301 16838 9331 16890
rect 9355 16838 9365 16890
rect 9365 16838 9411 16890
rect 9115 16836 9171 16838
rect 9195 16836 9251 16838
rect 9275 16836 9331 16838
rect 9355 16836 9411 16838
rect 9115 15802 9171 15804
rect 9195 15802 9251 15804
rect 9275 15802 9331 15804
rect 9355 15802 9411 15804
rect 9115 15750 9161 15802
rect 9161 15750 9171 15802
rect 9195 15750 9225 15802
rect 9225 15750 9237 15802
rect 9237 15750 9251 15802
rect 9275 15750 9289 15802
rect 9289 15750 9301 15802
rect 9301 15750 9331 15802
rect 9355 15750 9365 15802
rect 9365 15750 9411 15802
rect 9115 15748 9171 15750
rect 9195 15748 9251 15750
rect 9275 15748 9331 15750
rect 9355 15748 9411 15750
rect 10046 21528 10102 21584
rect 10046 20848 10102 20904
rect 10046 20032 10102 20088
rect 10046 19352 10102 19408
rect 10046 18572 10048 18592
rect 10048 18572 10100 18592
rect 10100 18572 10102 18592
rect 10046 18536 10102 18572
rect 10046 17720 10102 17776
rect 10046 17060 10102 17096
rect 10046 17040 10048 17060
rect 10048 17040 10100 17060
rect 10100 17040 10102 17060
rect 10046 16224 10102 16280
rect 10046 15544 10102 15600
rect 10046 14764 10048 14784
rect 10048 14764 10100 14784
rect 10100 14764 10102 14784
rect 10046 14728 10102 14764
rect 9115 14714 9171 14716
rect 9195 14714 9251 14716
rect 9275 14714 9331 14716
rect 9355 14714 9411 14716
rect 9115 14662 9161 14714
rect 9161 14662 9171 14714
rect 9195 14662 9225 14714
rect 9225 14662 9237 14714
rect 9237 14662 9251 14714
rect 9275 14662 9289 14714
rect 9289 14662 9301 14714
rect 9301 14662 9331 14714
rect 9355 14662 9365 14714
rect 9365 14662 9411 14714
rect 9115 14660 9171 14662
rect 9195 14660 9251 14662
rect 9275 14660 9331 14662
rect 9355 14660 9411 14662
rect 9115 13626 9171 13628
rect 9195 13626 9251 13628
rect 9275 13626 9331 13628
rect 9355 13626 9411 13628
rect 9115 13574 9161 13626
rect 9161 13574 9171 13626
rect 9195 13574 9225 13626
rect 9225 13574 9237 13626
rect 9237 13574 9251 13626
rect 9275 13574 9289 13626
rect 9289 13574 9301 13626
rect 9301 13574 9331 13626
rect 9355 13574 9365 13626
rect 9365 13574 9411 13626
rect 9115 13572 9171 13574
rect 9195 13572 9251 13574
rect 9275 13572 9331 13574
rect 9355 13572 9411 13574
rect 9115 12538 9171 12540
rect 9195 12538 9251 12540
rect 9275 12538 9331 12540
rect 9355 12538 9411 12540
rect 9115 12486 9161 12538
rect 9161 12486 9171 12538
rect 9195 12486 9225 12538
rect 9225 12486 9237 12538
rect 9237 12486 9251 12538
rect 9275 12486 9289 12538
rect 9289 12486 9301 12538
rect 9301 12486 9331 12538
rect 9355 12486 9365 12538
rect 9365 12486 9411 12538
rect 9115 12484 9171 12486
rect 9195 12484 9251 12486
rect 9275 12484 9331 12486
rect 9355 12484 9411 12486
rect 10046 13912 10102 13968
rect 10046 13232 10102 13288
rect 10046 12416 10102 12472
rect 10046 11736 10102 11792
rect 9115 11450 9171 11452
rect 9195 11450 9251 11452
rect 9275 11450 9331 11452
rect 9355 11450 9411 11452
rect 9115 11398 9161 11450
rect 9161 11398 9171 11450
rect 9195 11398 9225 11450
rect 9225 11398 9237 11450
rect 9237 11398 9251 11450
rect 9275 11398 9289 11450
rect 9289 11398 9301 11450
rect 9301 11398 9331 11450
rect 9355 11398 9365 11450
rect 9365 11398 9411 11450
rect 9115 11396 9171 11398
rect 9195 11396 9251 11398
rect 9275 11396 9331 11398
rect 9355 11396 9411 11398
rect 10046 10956 10048 10976
rect 10048 10956 10100 10976
rect 10100 10956 10102 10976
rect 10046 10920 10102 10956
rect 9115 10362 9171 10364
rect 9195 10362 9251 10364
rect 9275 10362 9331 10364
rect 9355 10362 9411 10364
rect 9115 10310 9161 10362
rect 9161 10310 9171 10362
rect 9195 10310 9225 10362
rect 9225 10310 9237 10362
rect 9237 10310 9251 10362
rect 9275 10310 9289 10362
rect 9289 10310 9301 10362
rect 9301 10310 9331 10362
rect 9355 10310 9365 10362
rect 9365 10310 9411 10362
rect 9115 10308 9171 10310
rect 9195 10308 9251 10310
rect 9275 10308 9331 10310
rect 9355 10308 9411 10310
rect 10046 10104 10102 10160
rect 10046 9444 10102 9480
rect 10046 9424 10048 9444
rect 10048 9424 10100 9444
rect 10100 9424 10102 9444
rect 9115 9274 9171 9276
rect 9195 9274 9251 9276
rect 9275 9274 9331 9276
rect 9355 9274 9411 9276
rect 9115 9222 9161 9274
rect 9161 9222 9171 9274
rect 9195 9222 9225 9274
rect 9225 9222 9237 9274
rect 9237 9222 9251 9274
rect 9275 9222 9289 9274
rect 9289 9222 9301 9274
rect 9301 9222 9331 9274
rect 9355 9222 9365 9274
rect 9365 9222 9411 9274
rect 9115 9220 9171 9222
rect 9195 9220 9251 9222
rect 9275 9220 9331 9222
rect 9355 9220 9411 9222
rect 10046 8608 10102 8664
rect 9115 8186 9171 8188
rect 9195 8186 9251 8188
rect 9275 8186 9331 8188
rect 9355 8186 9411 8188
rect 9115 8134 9161 8186
rect 9161 8134 9171 8186
rect 9195 8134 9225 8186
rect 9225 8134 9237 8186
rect 9237 8134 9251 8186
rect 9275 8134 9289 8186
rect 9289 8134 9301 8186
rect 9301 8134 9331 8186
rect 9355 8134 9365 8186
rect 9365 8134 9411 8186
rect 9115 8132 9171 8134
rect 9195 8132 9251 8134
rect 9275 8132 9331 8134
rect 9355 8132 9411 8134
rect 10046 7928 10102 7984
rect 7483 3290 7539 3292
rect 7563 3290 7619 3292
rect 7643 3290 7699 3292
rect 7723 3290 7779 3292
rect 7483 3238 7529 3290
rect 7529 3238 7539 3290
rect 7563 3238 7593 3290
rect 7593 3238 7605 3290
rect 7605 3238 7619 3290
rect 7643 3238 7657 3290
rect 7657 3238 7669 3290
rect 7669 3238 7699 3290
rect 7723 3238 7733 3290
rect 7733 3238 7779 3290
rect 7483 3236 7539 3238
rect 7563 3236 7619 3238
rect 7643 3236 7699 3238
rect 7723 3236 7779 3238
rect 5851 2746 5907 2748
rect 5931 2746 5987 2748
rect 6011 2746 6067 2748
rect 6091 2746 6147 2748
rect 5851 2694 5897 2746
rect 5897 2694 5907 2746
rect 5931 2694 5961 2746
rect 5961 2694 5973 2746
rect 5973 2694 5987 2746
rect 6011 2694 6025 2746
rect 6025 2694 6037 2746
rect 6037 2694 6067 2746
rect 6091 2694 6101 2746
rect 6101 2694 6147 2746
rect 5851 2692 5907 2694
rect 5931 2692 5987 2694
rect 6011 2692 6067 2694
rect 6091 2692 6147 2694
rect 9115 7098 9171 7100
rect 9195 7098 9251 7100
rect 9275 7098 9331 7100
rect 9355 7098 9411 7100
rect 9115 7046 9161 7098
rect 9161 7046 9171 7098
rect 9195 7046 9225 7098
rect 9225 7046 9237 7098
rect 9237 7046 9251 7098
rect 9275 7046 9289 7098
rect 9289 7046 9301 7098
rect 9301 7046 9331 7098
rect 9355 7046 9365 7098
rect 9365 7046 9411 7098
rect 9115 7044 9171 7046
rect 9195 7044 9251 7046
rect 9275 7044 9331 7046
rect 9355 7044 9411 7046
rect 9115 6010 9171 6012
rect 9195 6010 9251 6012
rect 9275 6010 9331 6012
rect 9355 6010 9411 6012
rect 9115 5958 9161 6010
rect 9161 5958 9171 6010
rect 9195 5958 9225 6010
rect 9225 5958 9237 6010
rect 9237 5958 9251 6010
rect 9275 5958 9289 6010
rect 9289 5958 9301 6010
rect 9301 5958 9331 6010
rect 9355 5958 9365 6010
rect 9365 5958 9411 6010
rect 9115 5956 9171 5958
rect 9195 5956 9251 5958
rect 9275 5956 9331 5958
rect 9355 5956 9411 5958
rect 10046 7148 10048 7168
rect 10048 7148 10100 7168
rect 10100 7148 10102 7168
rect 10046 7112 10102 7148
rect 9115 4922 9171 4924
rect 9195 4922 9251 4924
rect 9275 4922 9331 4924
rect 9355 4922 9411 4924
rect 9115 4870 9161 4922
rect 9161 4870 9171 4922
rect 9195 4870 9225 4922
rect 9225 4870 9237 4922
rect 9237 4870 9251 4922
rect 9275 4870 9289 4922
rect 9289 4870 9301 4922
rect 9301 4870 9331 4922
rect 9355 4870 9365 4922
rect 9365 4870 9411 4922
rect 9115 4868 9171 4870
rect 9195 4868 9251 4870
rect 9275 4868 9331 4870
rect 9355 4868 9411 4870
rect 10046 6296 10102 6352
rect 10046 5616 10102 5672
rect 10046 4800 10102 4856
rect 9115 3834 9171 3836
rect 9195 3834 9251 3836
rect 9275 3834 9331 3836
rect 9355 3834 9411 3836
rect 9115 3782 9161 3834
rect 9161 3782 9171 3834
rect 9195 3782 9225 3834
rect 9225 3782 9237 3834
rect 9237 3782 9251 3834
rect 9275 3782 9289 3834
rect 9289 3782 9301 3834
rect 9301 3782 9331 3834
rect 9355 3782 9365 3834
rect 9365 3782 9411 3834
rect 9115 3780 9171 3782
rect 9195 3780 9251 3782
rect 9275 3780 9331 3782
rect 9355 3780 9411 3782
rect 9115 2746 9171 2748
rect 9195 2746 9251 2748
rect 9275 2746 9331 2748
rect 9355 2746 9411 2748
rect 9115 2694 9161 2746
rect 9161 2694 9171 2746
rect 9195 2694 9225 2746
rect 9225 2694 9237 2746
rect 9237 2694 9251 2746
rect 9275 2694 9289 2746
rect 9289 2694 9301 2746
rect 9301 2694 9331 2746
rect 9355 2694 9365 2746
rect 9365 2694 9411 2746
rect 9115 2692 9171 2694
rect 9195 2692 9251 2694
rect 9275 2692 9331 2694
rect 9355 2692 9411 2694
rect 4219 2202 4275 2204
rect 4299 2202 4355 2204
rect 4379 2202 4435 2204
rect 4459 2202 4515 2204
rect 4219 2150 4265 2202
rect 4265 2150 4275 2202
rect 4299 2150 4329 2202
rect 4329 2150 4341 2202
rect 4341 2150 4355 2202
rect 4379 2150 4393 2202
rect 4393 2150 4405 2202
rect 4405 2150 4435 2202
rect 4459 2150 4469 2202
rect 4469 2150 4515 2202
rect 4219 2148 4275 2150
rect 4299 2148 4355 2150
rect 4379 2148 4435 2150
rect 4459 2148 4515 2150
rect 3974 1808 4030 1864
rect 3606 992 3662 1048
rect 2778 584 2834 640
rect 7483 2202 7539 2204
rect 7563 2202 7619 2204
rect 7643 2202 7699 2204
rect 7723 2202 7779 2204
rect 7483 2150 7529 2202
rect 7529 2150 7539 2202
rect 7563 2150 7593 2202
rect 7593 2150 7605 2202
rect 7605 2150 7619 2202
rect 7643 2150 7657 2202
rect 7657 2150 7669 2202
rect 7669 2150 7699 2202
rect 7723 2150 7733 2202
rect 7733 2150 7779 2202
rect 7483 2148 7539 2150
rect 7563 2148 7619 2150
rect 7643 2148 7699 2150
rect 7723 2148 7779 2150
rect 2778 176 2834 232
rect 10046 4120 10102 4176
rect 10046 3340 10048 3360
rect 10048 3340 10100 3360
rect 10100 3340 10102 3360
rect 10046 3304 10102 3340
rect 10046 2488 10102 2544
rect 9494 1808 9550 1864
rect 10046 992 10102 1048
rect 9310 312 9366 368
<< metal3 >>
rect 0 79658 800 79688
rect 2957 79658 3023 79661
rect 0 79656 3023 79658
rect 0 79600 2962 79656
rect 3018 79600 3023 79656
rect 0 79598 3023 79600
rect 0 79568 800 79598
rect 2957 79595 3023 79598
rect 11200 79432 12000 79552
rect 0 79250 800 79280
rect 3877 79250 3943 79253
rect 0 79248 3943 79250
rect 0 79192 3882 79248
rect 3938 79192 3943 79248
rect 0 79190 3943 79192
rect 0 79160 800 79190
rect 3877 79187 3943 79190
rect 0 78842 800 78872
rect 3049 78842 3115 78845
rect 0 78840 3115 78842
rect 0 78784 3054 78840
rect 3110 78784 3115 78840
rect 0 78782 3115 78784
rect 0 78752 800 78782
rect 3049 78779 3115 78782
rect 10133 78706 10199 78709
rect 11200 78706 12000 78736
rect 10133 78704 12000 78706
rect 10133 78648 10138 78704
rect 10194 78648 12000 78704
rect 10133 78646 12000 78648
rect 10133 78643 10199 78646
rect 11200 78616 12000 78646
rect 0 78434 800 78464
rect 3325 78434 3391 78437
rect 0 78432 3391 78434
rect 0 78376 3330 78432
rect 3386 78376 3391 78432
rect 0 78374 3391 78376
rect 0 78344 800 78374
rect 3325 78371 3391 78374
rect 0 78026 800 78056
rect 4061 78026 4127 78029
rect 0 78024 4127 78026
rect 0 77968 4066 78024
rect 4122 77968 4127 78024
rect 0 77966 4127 77968
rect 0 77936 800 77966
rect 4061 77963 4127 77966
rect 10961 78026 11027 78029
rect 11200 78026 12000 78056
rect 10961 78024 12000 78026
rect 10961 77968 10966 78024
rect 11022 77968 12000 78024
rect 10961 77966 12000 77968
rect 10961 77963 11027 77966
rect 11200 77936 12000 77966
rect 2576 77824 2896 77825
rect 2576 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2576 77759 2896 77760
rect 5839 77824 6159 77825
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 77759 6159 77760
rect 9103 77824 9423 77825
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 77759 9423 77760
rect 0 77618 800 77648
rect 3969 77618 4035 77621
rect 0 77616 4035 77618
rect 0 77560 3974 77616
rect 4030 77560 4035 77616
rect 0 77558 4035 77560
rect 0 77528 800 77558
rect 3969 77555 4035 77558
rect 4207 77280 4527 77281
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 77215 4527 77216
rect 7471 77280 7791 77281
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 77215 7791 77216
rect 9397 77210 9463 77213
rect 11200 77210 12000 77240
rect 9397 77208 12000 77210
rect 9397 77152 9402 77208
rect 9458 77152 12000 77208
rect 9397 77150 12000 77152
rect 9397 77147 9463 77150
rect 11200 77120 12000 77150
rect 0 77074 800 77104
rect 2497 77074 2563 77077
rect 0 77072 2563 77074
rect 0 77016 2502 77072
rect 2558 77016 2563 77072
rect 0 77014 2563 77016
rect 0 76984 800 77014
rect 2497 77011 2563 77014
rect 2773 76938 2839 76941
rect 1396 76936 2839 76938
rect 1396 76880 2778 76936
rect 2834 76880 2839 76936
rect 1396 76878 2839 76880
rect 0 76666 800 76696
rect 1396 76666 1456 76878
rect 2773 76875 2839 76878
rect 2576 76736 2896 76737
rect 2576 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2576 76671 2896 76672
rect 5839 76736 6159 76737
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 76671 6159 76672
rect 9103 76736 9423 76737
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 76671 9423 76672
rect 0 76606 1456 76666
rect 0 76576 800 76606
rect 10133 76530 10199 76533
rect 11200 76530 12000 76560
rect 10133 76528 12000 76530
rect 10133 76472 10138 76528
rect 10194 76472 12000 76528
rect 10133 76470 12000 76472
rect 10133 76467 10199 76470
rect 11200 76440 12000 76470
rect 0 76258 800 76288
rect 2037 76258 2103 76261
rect 0 76256 2103 76258
rect 0 76200 2042 76256
rect 2098 76200 2103 76256
rect 0 76198 2103 76200
rect 0 76168 800 76198
rect 2037 76195 2103 76198
rect 4207 76192 4527 76193
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 76127 4527 76128
rect 7471 76192 7791 76193
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 76127 7791 76128
rect 0 75850 800 75880
rect 2957 75850 3023 75853
rect 0 75848 3023 75850
rect 0 75792 2962 75848
rect 3018 75792 3023 75848
rect 0 75790 3023 75792
rect 0 75760 800 75790
rect 2957 75787 3023 75790
rect 10225 75714 10291 75717
rect 11200 75714 12000 75744
rect 10225 75712 12000 75714
rect 10225 75656 10230 75712
rect 10286 75656 12000 75712
rect 10225 75654 12000 75656
rect 10225 75651 10291 75654
rect 2576 75648 2896 75649
rect 2576 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2576 75583 2896 75584
rect 5839 75648 6159 75649
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 75583 6159 75584
rect 9103 75648 9423 75649
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 11200 75624 12000 75654
rect 9103 75583 9423 75584
rect 0 75442 800 75472
rect 1393 75442 1459 75445
rect 0 75440 1459 75442
rect 0 75384 1398 75440
rect 1454 75384 1459 75440
rect 0 75382 1459 75384
rect 0 75352 800 75382
rect 1393 75379 1459 75382
rect 4207 75104 4527 75105
rect 0 75034 800 75064
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 75039 4527 75040
rect 7471 75104 7791 75105
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 75039 7791 75040
rect 3969 75034 4035 75037
rect 0 75032 4035 75034
rect 0 74976 3974 75032
rect 4030 74976 4035 75032
rect 0 74974 4035 74976
rect 0 74944 800 74974
rect 3969 74971 4035 74974
rect 10133 74898 10199 74901
rect 11200 74898 12000 74928
rect 10133 74896 12000 74898
rect 10133 74840 10138 74896
rect 10194 74840 12000 74896
rect 10133 74838 12000 74840
rect 10133 74835 10199 74838
rect 11200 74808 12000 74838
rect 2576 74560 2896 74561
rect 0 74490 800 74520
rect 2576 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2576 74495 2896 74496
rect 5839 74560 6159 74561
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 74495 6159 74496
rect 9103 74560 9423 74561
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 74495 9423 74496
rect 0 74430 1456 74490
rect 0 74400 800 74430
rect 1396 74354 1456 74430
rect 3601 74354 3667 74357
rect 1396 74352 3667 74354
rect 1396 74296 3606 74352
rect 3662 74296 3667 74352
rect 1396 74294 3667 74296
rect 3601 74291 3667 74294
rect 10133 74218 10199 74221
rect 11200 74218 12000 74248
rect 10133 74216 12000 74218
rect 10133 74160 10138 74216
rect 10194 74160 12000 74216
rect 10133 74158 12000 74160
rect 10133 74155 10199 74158
rect 11200 74128 12000 74158
rect 0 74082 800 74112
rect 1301 74082 1367 74085
rect 0 74080 1367 74082
rect 0 74024 1306 74080
rect 1362 74024 1367 74080
rect 0 74022 1367 74024
rect 0 73992 800 74022
rect 1301 74019 1367 74022
rect 4207 74016 4527 74017
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 73951 4527 73952
rect 7471 74016 7791 74017
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 73951 7791 73952
rect 0 73674 800 73704
rect 1393 73674 1459 73677
rect 0 73672 1459 73674
rect 0 73616 1398 73672
rect 1454 73616 1459 73672
rect 0 73614 1459 73616
rect 0 73584 800 73614
rect 1393 73611 1459 73614
rect 2576 73472 2896 73473
rect 2576 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2576 73407 2896 73408
rect 5839 73472 6159 73473
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 73407 6159 73408
rect 9103 73472 9423 73473
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 73407 9423 73408
rect 10133 73402 10199 73405
rect 11200 73402 12000 73432
rect 10133 73400 12000 73402
rect 10133 73344 10138 73400
rect 10194 73344 12000 73400
rect 10133 73342 12000 73344
rect 10133 73339 10199 73342
rect 11200 73312 12000 73342
rect 0 73266 800 73296
rect 2957 73266 3023 73269
rect 0 73264 3023 73266
rect 0 73208 2962 73264
rect 3018 73208 3023 73264
rect 0 73206 3023 73208
rect 0 73176 800 73206
rect 2957 73203 3023 73206
rect 4207 72928 4527 72929
rect 0 72858 800 72888
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 72863 4527 72864
rect 7471 72928 7791 72929
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 72863 7791 72864
rect 2221 72858 2287 72861
rect 0 72856 2287 72858
rect 0 72800 2226 72856
rect 2282 72800 2287 72856
rect 0 72798 2287 72800
rect 0 72768 800 72798
rect 2221 72795 2287 72798
rect 10133 72722 10199 72725
rect 11200 72722 12000 72752
rect 10133 72720 12000 72722
rect 10133 72664 10138 72720
rect 10194 72664 12000 72720
rect 10133 72662 12000 72664
rect 10133 72659 10199 72662
rect 11200 72632 12000 72662
rect 0 72450 800 72480
rect 1393 72450 1459 72453
rect 0 72448 1459 72450
rect 0 72392 1398 72448
rect 1454 72392 1459 72448
rect 0 72390 1459 72392
rect 0 72360 800 72390
rect 1393 72387 1459 72390
rect 2576 72384 2896 72385
rect 2576 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2576 72319 2896 72320
rect 5839 72384 6159 72385
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 72319 6159 72320
rect 9103 72384 9423 72385
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 72319 9423 72320
rect 1761 72178 1827 72181
rect 2129 72178 2195 72181
rect 1761 72176 2195 72178
rect 1761 72120 1766 72176
rect 1822 72120 2134 72176
rect 2190 72120 2195 72176
rect 1761 72118 2195 72120
rect 1761 72115 1827 72118
rect 2129 72115 2195 72118
rect 0 71906 800 71936
rect 1301 71906 1367 71909
rect 0 71904 1367 71906
rect 0 71848 1306 71904
rect 1362 71848 1367 71904
rect 0 71846 1367 71848
rect 0 71816 800 71846
rect 1301 71843 1367 71846
rect 10133 71906 10199 71909
rect 11200 71906 12000 71936
rect 10133 71904 12000 71906
rect 10133 71848 10138 71904
rect 10194 71848 12000 71904
rect 10133 71846 12000 71848
rect 10133 71843 10199 71846
rect 4207 71840 4527 71841
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 71775 4527 71776
rect 7471 71840 7791 71841
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 11200 71816 12000 71846
rect 7471 71775 7791 71776
rect 0 71498 800 71528
rect 1301 71498 1367 71501
rect 0 71496 1367 71498
rect 0 71440 1306 71496
rect 1362 71440 1367 71496
rect 0 71438 1367 71440
rect 0 71408 800 71438
rect 1301 71435 1367 71438
rect 2576 71296 2896 71297
rect 2576 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2576 71231 2896 71232
rect 5839 71296 6159 71297
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 71231 6159 71232
rect 9103 71296 9423 71297
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 71231 9423 71232
rect 0 71090 800 71120
rect 1393 71090 1459 71093
rect 0 71088 1459 71090
rect 0 71032 1398 71088
rect 1454 71032 1459 71088
rect 0 71030 1459 71032
rect 0 71000 800 71030
rect 1393 71027 1459 71030
rect 10133 71090 10199 71093
rect 11200 71090 12000 71120
rect 10133 71088 12000 71090
rect 10133 71032 10138 71088
rect 10194 71032 12000 71088
rect 10133 71030 12000 71032
rect 10133 71027 10199 71030
rect 11200 71000 12000 71030
rect 4207 70752 4527 70753
rect 0 70682 800 70712
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 70687 4527 70688
rect 7471 70752 7791 70753
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 70687 7791 70688
rect 2773 70682 2839 70685
rect 0 70680 2839 70682
rect 0 70624 2778 70680
rect 2834 70624 2839 70680
rect 0 70622 2839 70624
rect 0 70592 800 70622
rect 2773 70619 2839 70622
rect 10133 70410 10199 70413
rect 11200 70410 12000 70440
rect 10133 70408 12000 70410
rect 10133 70352 10138 70408
rect 10194 70352 12000 70408
rect 10133 70350 12000 70352
rect 10133 70347 10199 70350
rect 11200 70320 12000 70350
rect 0 70274 800 70304
rect 1301 70274 1367 70277
rect 0 70272 1367 70274
rect 0 70216 1306 70272
rect 1362 70216 1367 70272
rect 0 70214 1367 70216
rect 0 70184 800 70214
rect 1301 70211 1367 70214
rect 2576 70208 2896 70209
rect 2576 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2576 70143 2896 70144
rect 5839 70208 6159 70209
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 70143 6159 70144
rect 9103 70208 9423 70209
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 70143 9423 70144
rect 0 69866 800 69896
rect 3509 69866 3575 69869
rect 0 69864 3575 69866
rect 0 69808 3514 69864
rect 3570 69808 3575 69864
rect 0 69806 3575 69808
rect 0 69776 800 69806
rect 3509 69803 3575 69806
rect 1577 69730 1643 69733
rect 2405 69730 2471 69733
rect 1577 69728 2471 69730
rect 1577 69672 1582 69728
rect 1638 69672 2410 69728
rect 2466 69672 2471 69728
rect 1577 69670 2471 69672
rect 1577 69667 1643 69670
rect 2405 69667 2471 69670
rect 4207 69664 4527 69665
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 69599 4527 69600
rect 7471 69664 7791 69665
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 69599 7791 69600
rect 10133 69594 10199 69597
rect 11200 69594 12000 69624
rect 10133 69592 12000 69594
rect 10133 69536 10138 69592
rect 10194 69536 12000 69592
rect 10133 69534 12000 69536
rect 10133 69531 10199 69534
rect 11200 69504 12000 69534
rect 1761 69458 1827 69461
rect 5717 69458 5783 69461
rect 1761 69456 5783 69458
rect 1761 69400 1766 69456
rect 1822 69400 5722 69456
rect 5778 69400 5783 69456
rect 1761 69398 5783 69400
rect 1761 69395 1827 69398
rect 5717 69395 5783 69398
rect 0 69322 800 69352
rect 3969 69322 4035 69325
rect 0 69320 4035 69322
rect 0 69264 3974 69320
rect 4030 69264 4035 69320
rect 0 69262 4035 69264
rect 0 69232 800 69262
rect 3969 69259 4035 69262
rect 2576 69120 2896 69121
rect 2576 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 2576 69055 2896 69056
rect 5839 69120 6159 69121
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 69055 6159 69056
rect 9103 69120 9423 69121
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 69055 9423 69056
rect 1158 68988 1164 69052
rect 1228 69050 1234 69052
rect 1485 69050 1551 69053
rect 1228 69048 1551 69050
rect 1228 68992 1490 69048
rect 1546 68992 1551 69048
rect 1228 68990 1551 68992
rect 1228 68988 1234 68990
rect 1485 68987 1551 68990
rect 0 68914 800 68944
rect 4153 68914 4219 68917
rect 0 68912 4219 68914
rect 0 68856 4158 68912
rect 4214 68856 4219 68912
rect 0 68854 4219 68856
rect 0 68824 800 68854
rect 4153 68851 4219 68854
rect 10133 68914 10199 68917
rect 11200 68914 12000 68944
rect 10133 68912 12000 68914
rect 10133 68856 10138 68912
rect 10194 68856 12000 68912
rect 10133 68854 12000 68856
rect 10133 68851 10199 68854
rect 11200 68824 12000 68854
rect 4207 68576 4527 68577
rect 0 68506 800 68536
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 68511 4527 68512
rect 7471 68576 7791 68577
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 68511 7791 68512
rect 3969 68506 4035 68509
rect 0 68504 4035 68506
rect 0 68448 3974 68504
rect 4030 68448 4035 68504
rect 0 68446 4035 68448
rect 0 68416 800 68446
rect 3969 68443 4035 68446
rect 3417 68234 3483 68237
rect 1350 68232 3483 68234
rect 1350 68176 3422 68232
rect 3478 68176 3483 68232
rect 1350 68174 3483 68176
rect 0 68098 800 68128
rect 1350 68098 1410 68174
rect 3417 68171 3483 68174
rect 0 68038 1410 68098
rect 10133 68098 10199 68101
rect 11200 68098 12000 68128
rect 10133 68096 12000 68098
rect 10133 68040 10138 68096
rect 10194 68040 12000 68096
rect 10133 68038 12000 68040
rect 0 68008 800 68038
rect 10133 68035 10199 68038
rect 2576 68032 2896 68033
rect 2576 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2576 67967 2896 67968
rect 5839 68032 6159 68033
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 67967 6159 67968
rect 9103 68032 9423 68033
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 11200 68008 12000 68038
rect 9103 67967 9423 67968
rect 0 67690 800 67720
rect 1301 67690 1367 67693
rect 0 67688 1367 67690
rect 0 67632 1306 67688
rect 1362 67632 1367 67688
rect 0 67630 1367 67632
rect 0 67600 800 67630
rect 1301 67627 1367 67630
rect 4207 67488 4527 67489
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 67423 4527 67424
rect 7471 67488 7791 67489
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 67423 7791 67424
rect 0 67282 800 67312
rect 1393 67282 1459 67285
rect 0 67280 1459 67282
rect 0 67224 1398 67280
rect 1454 67224 1459 67280
rect 0 67222 1459 67224
rect 0 67192 800 67222
rect 1393 67219 1459 67222
rect 10133 67282 10199 67285
rect 11200 67282 12000 67312
rect 10133 67280 12000 67282
rect 10133 67224 10138 67280
rect 10194 67224 12000 67280
rect 10133 67222 12000 67224
rect 10133 67219 10199 67222
rect 11200 67192 12000 67222
rect 2576 66944 2896 66945
rect 0 66874 800 66904
rect 2576 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2576 66879 2896 66880
rect 5839 66944 6159 66945
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 66879 6159 66880
rect 9103 66944 9423 66945
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 66879 9423 66880
rect 0 66814 1410 66874
rect 0 66784 800 66814
rect 1350 66738 1410 66814
rect 2957 66738 3023 66741
rect 1350 66736 3023 66738
rect 1350 66680 2962 66736
rect 3018 66680 3023 66736
rect 1350 66678 3023 66680
rect 2957 66675 3023 66678
rect 10133 66602 10199 66605
rect 11200 66602 12000 66632
rect 10133 66600 12000 66602
rect 10133 66544 10138 66600
rect 10194 66544 12000 66600
rect 10133 66542 12000 66544
rect 10133 66539 10199 66542
rect 11200 66512 12000 66542
rect 4207 66400 4527 66401
rect 0 66330 800 66360
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 66335 4527 66336
rect 7471 66400 7791 66401
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 66335 7791 66336
rect 2313 66330 2379 66333
rect 0 66328 2379 66330
rect 0 66272 2318 66328
rect 2374 66272 2379 66328
rect 0 66270 2379 66272
rect 0 66240 800 66270
rect 2313 66267 2379 66270
rect 0 65922 800 65952
rect 1393 65922 1459 65925
rect 0 65920 1459 65922
rect 0 65864 1398 65920
rect 1454 65864 1459 65920
rect 0 65862 1459 65864
rect 0 65832 800 65862
rect 1393 65859 1459 65862
rect 2576 65856 2896 65857
rect 2576 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2576 65791 2896 65792
rect 5839 65856 6159 65857
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 65791 6159 65792
rect 9103 65856 9423 65857
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 65791 9423 65792
rect 10133 65786 10199 65789
rect 11200 65786 12000 65816
rect 10133 65784 12000 65786
rect 10133 65728 10138 65784
rect 10194 65728 12000 65784
rect 10133 65726 12000 65728
rect 10133 65723 10199 65726
rect 11200 65696 12000 65726
rect 0 65514 800 65544
rect 1485 65514 1551 65517
rect 0 65512 1551 65514
rect 0 65456 1490 65512
rect 1546 65456 1551 65512
rect 0 65454 1551 65456
rect 0 65424 800 65454
rect 1485 65451 1551 65454
rect 4207 65312 4527 65313
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 65247 4527 65248
rect 7471 65312 7791 65313
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 65247 7791 65248
rect 0 65106 800 65136
rect 3049 65106 3115 65109
rect 0 65104 3115 65106
rect 0 65048 3054 65104
rect 3110 65048 3115 65104
rect 0 65046 3115 65048
rect 0 65016 800 65046
rect 3049 65043 3115 65046
rect 10133 65106 10199 65109
rect 11200 65106 12000 65136
rect 10133 65104 12000 65106
rect 10133 65048 10138 65104
rect 10194 65048 12000 65104
rect 10133 65046 12000 65048
rect 10133 65043 10199 65046
rect 11200 65016 12000 65046
rect 2313 64834 2379 64837
rect 1166 64832 2379 64834
rect 1166 64776 2318 64832
rect 2374 64776 2379 64832
rect 1166 64774 2379 64776
rect 0 64698 800 64728
rect 1166 64698 1226 64774
rect 2313 64771 2379 64774
rect 2576 64768 2896 64769
rect 2576 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2576 64703 2896 64704
rect 5839 64768 6159 64769
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 64703 6159 64704
rect 9103 64768 9423 64769
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 64703 9423 64704
rect 0 64638 1226 64698
rect 0 64608 800 64638
rect 0 64290 800 64320
rect 1485 64290 1551 64293
rect 0 64288 1551 64290
rect 0 64232 1490 64288
rect 1546 64232 1551 64288
rect 0 64230 1551 64232
rect 0 64200 800 64230
rect 1485 64227 1551 64230
rect 10133 64290 10199 64293
rect 11200 64290 12000 64320
rect 10133 64288 12000 64290
rect 10133 64232 10138 64288
rect 10194 64232 12000 64288
rect 10133 64230 12000 64232
rect 10133 64227 10199 64230
rect 4207 64224 4527 64225
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 64159 4527 64160
rect 7471 64224 7791 64225
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 11200 64200 12000 64230
rect 7471 64159 7791 64160
rect 3877 63882 3943 63885
rect 1350 63880 3943 63882
rect 1350 63824 3882 63880
rect 3938 63824 3943 63880
rect 1350 63822 3943 63824
rect 0 63746 800 63776
rect 1350 63746 1410 63822
rect 3877 63819 3943 63822
rect 0 63686 1410 63746
rect 0 63656 800 63686
rect 2576 63680 2896 63681
rect 2576 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2576 63615 2896 63616
rect 5839 63680 6159 63681
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 63615 6159 63616
rect 9103 63680 9423 63681
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 63615 9423 63616
rect 2865 63474 2931 63477
rect 4061 63474 4127 63477
rect 2865 63472 4127 63474
rect 2865 63416 2870 63472
rect 2926 63416 4066 63472
rect 4122 63416 4127 63472
rect 2865 63414 4127 63416
rect 2865 63411 2931 63414
rect 4061 63411 4127 63414
rect 10133 63474 10199 63477
rect 11200 63474 12000 63504
rect 10133 63472 12000 63474
rect 10133 63416 10138 63472
rect 10194 63416 12000 63472
rect 10133 63414 12000 63416
rect 10133 63411 10199 63414
rect 11200 63384 12000 63414
rect 0 63338 800 63368
rect 3141 63338 3207 63341
rect 0 63336 3207 63338
rect 0 63280 3146 63336
rect 3202 63280 3207 63336
rect 0 63278 3207 63280
rect 0 63248 800 63278
rect 3141 63275 3207 63278
rect 2865 63202 2931 63205
rect 4061 63202 4127 63205
rect 2865 63200 4127 63202
rect 2865 63144 2870 63200
rect 2926 63144 4066 63200
rect 4122 63144 4127 63200
rect 2865 63142 4127 63144
rect 2865 63139 2931 63142
rect 4061 63139 4127 63142
rect 4207 63136 4527 63137
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 63071 4527 63072
rect 7471 63136 7791 63137
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 63071 7791 63072
rect 0 62930 800 62960
rect 3969 62930 4035 62933
rect 0 62928 4035 62930
rect 0 62872 3974 62928
rect 4030 62872 4035 62928
rect 0 62870 4035 62872
rect 0 62840 800 62870
rect 3969 62867 4035 62870
rect 10133 62794 10199 62797
rect 11200 62794 12000 62824
rect 10133 62792 12000 62794
rect 10133 62736 10138 62792
rect 10194 62736 12000 62792
rect 10133 62734 12000 62736
rect 10133 62731 10199 62734
rect 11200 62704 12000 62734
rect 2576 62592 2896 62593
rect 0 62522 800 62552
rect 2576 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2576 62527 2896 62528
rect 5839 62592 6159 62593
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 62527 6159 62528
rect 9103 62592 9423 62593
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 62527 9423 62528
rect 1393 62522 1459 62525
rect 0 62520 1459 62522
rect 0 62464 1398 62520
rect 1454 62464 1459 62520
rect 0 62462 1459 62464
rect 0 62432 800 62462
rect 1393 62459 1459 62462
rect 0 62114 800 62144
rect 2221 62114 2287 62117
rect 0 62112 2287 62114
rect 0 62056 2226 62112
rect 2282 62056 2287 62112
rect 0 62054 2287 62056
rect 0 62024 800 62054
rect 2221 62051 2287 62054
rect 4207 62048 4527 62049
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 61983 4527 61984
rect 7471 62048 7791 62049
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 61983 7791 61984
rect 2037 61978 2103 61981
rect 2221 61978 2287 61981
rect 2037 61976 2287 61978
rect 2037 61920 2042 61976
rect 2098 61920 2226 61976
rect 2282 61920 2287 61976
rect 2037 61918 2287 61920
rect 2037 61915 2103 61918
rect 2221 61915 2287 61918
rect 10133 61978 10199 61981
rect 11200 61978 12000 62008
rect 10133 61976 12000 61978
rect 10133 61920 10138 61976
rect 10194 61920 12000 61976
rect 10133 61918 12000 61920
rect 10133 61915 10199 61918
rect 11200 61888 12000 61918
rect 0 61706 800 61736
rect 1485 61706 1551 61709
rect 0 61704 1551 61706
rect 0 61648 1490 61704
rect 1546 61648 1551 61704
rect 0 61646 1551 61648
rect 0 61616 800 61646
rect 1485 61643 1551 61646
rect 2576 61504 2896 61505
rect 2576 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2576 61439 2896 61440
rect 5839 61504 6159 61505
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 61439 6159 61440
rect 9103 61504 9423 61505
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 61439 9423 61440
rect 10133 61298 10199 61301
rect 11200 61298 12000 61328
rect 10133 61296 12000 61298
rect 10133 61240 10138 61296
rect 10194 61240 12000 61296
rect 10133 61238 12000 61240
rect 10133 61235 10199 61238
rect 11200 61208 12000 61238
rect 0 61162 800 61192
rect 3969 61162 4035 61165
rect 0 61160 4035 61162
rect 0 61104 3974 61160
rect 4030 61104 4035 61160
rect 0 61102 4035 61104
rect 0 61072 800 61102
rect 3969 61099 4035 61102
rect 4207 60960 4527 60961
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 60895 4527 60896
rect 7471 60960 7791 60961
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 60895 7791 60896
rect 0 60754 800 60784
rect 2957 60754 3023 60757
rect 0 60752 3023 60754
rect 0 60696 2962 60752
rect 3018 60696 3023 60752
rect 0 60694 3023 60696
rect 0 60664 800 60694
rect 2957 60691 3023 60694
rect 3325 60754 3391 60757
rect 3877 60754 3943 60757
rect 3325 60752 3943 60754
rect 3325 60696 3330 60752
rect 3386 60696 3882 60752
rect 3938 60696 3943 60752
rect 3325 60694 3943 60696
rect 3325 60691 3391 60694
rect 3877 60691 3943 60694
rect 5533 60754 5599 60757
rect 5533 60752 5642 60754
rect 5533 60696 5538 60752
rect 5594 60696 5642 60752
rect 5533 60691 5642 60696
rect 2773 60618 2839 60621
rect 1350 60616 2839 60618
rect 1350 60560 2778 60616
rect 2834 60560 2839 60616
rect 1350 60558 2839 60560
rect 5582 60618 5642 60691
rect 6177 60618 6243 60621
rect 5582 60616 6243 60618
rect 5582 60560 6182 60616
rect 6238 60560 6243 60616
rect 5582 60558 6243 60560
rect 0 60346 800 60376
rect 1350 60346 1410 60558
rect 2773 60555 2839 60558
rect 6177 60555 6243 60558
rect 10133 60482 10199 60485
rect 11200 60482 12000 60512
rect 10133 60480 12000 60482
rect 10133 60424 10138 60480
rect 10194 60424 12000 60480
rect 10133 60422 12000 60424
rect 10133 60419 10199 60422
rect 2576 60416 2896 60417
rect 2576 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2576 60351 2896 60352
rect 5839 60416 6159 60417
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 60351 6159 60352
rect 9103 60416 9423 60417
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 11200 60392 12000 60422
rect 9103 60351 9423 60352
rect 0 60286 1410 60346
rect 0 60256 800 60286
rect 0 59938 800 59968
rect 1485 59938 1551 59941
rect 0 59936 1551 59938
rect 0 59880 1490 59936
rect 1546 59880 1551 59936
rect 0 59878 1551 59880
rect 0 59848 800 59878
rect 1485 59875 1551 59878
rect 4207 59872 4527 59873
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 59807 4527 59808
rect 7471 59872 7791 59873
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 59807 7791 59808
rect 10133 59666 10199 59669
rect 11200 59666 12000 59696
rect 10133 59664 12000 59666
rect 10133 59608 10138 59664
rect 10194 59608 12000 59664
rect 10133 59606 12000 59608
rect 10133 59603 10199 59606
rect 11200 59576 12000 59606
rect 0 59530 800 59560
rect 1393 59530 1459 59533
rect 0 59528 1459 59530
rect 0 59472 1398 59528
rect 1454 59472 1459 59528
rect 0 59470 1459 59472
rect 0 59440 800 59470
rect 1393 59467 1459 59470
rect 2576 59328 2896 59329
rect 2576 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2576 59263 2896 59264
rect 5839 59328 6159 59329
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 59263 6159 59264
rect 9103 59328 9423 59329
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 59263 9423 59264
rect 0 59122 800 59152
rect 1301 59122 1367 59125
rect 0 59120 1367 59122
rect 0 59064 1306 59120
rect 1362 59064 1367 59120
rect 0 59062 1367 59064
rect 0 59032 800 59062
rect 1301 59059 1367 59062
rect 10133 58986 10199 58989
rect 11200 58986 12000 59016
rect 10133 58984 12000 58986
rect 10133 58928 10138 58984
rect 10194 58928 12000 58984
rect 10133 58926 12000 58928
rect 10133 58923 10199 58926
rect 11200 58896 12000 58926
rect 841 58850 907 58853
rect 798 58848 907 58850
rect 798 58792 846 58848
rect 902 58792 907 58848
rect 798 58787 907 58792
rect 798 58608 858 58787
rect 4207 58784 4527 58785
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 58719 4527 58720
rect 7471 58784 7791 58785
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 58719 7791 58720
rect 0 58518 858 58608
rect 0 58488 800 58518
rect 2576 58240 2896 58241
rect 0 58170 800 58200
rect 2576 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2576 58175 2896 58176
rect 5839 58240 6159 58241
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 58175 6159 58176
rect 9103 58240 9423 58241
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 58175 9423 58176
rect 1485 58170 1551 58173
rect 0 58168 1551 58170
rect 0 58112 1490 58168
rect 1546 58112 1551 58168
rect 0 58110 1551 58112
rect 0 58080 800 58110
rect 1485 58107 1551 58110
rect 10133 58170 10199 58173
rect 11200 58170 12000 58200
rect 10133 58168 12000 58170
rect 10133 58112 10138 58168
rect 10194 58112 12000 58168
rect 10133 58110 12000 58112
rect 10133 58107 10199 58110
rect 11200 58080 12000 58110
rect 1301 57898 1367 57901
rect 1853 57898 1919 57901
rect 1301 57896 1919 57898
rect 1301 57840 1306 57896
rect 1362 57840 1858 57896
rect 1914 57840 1919 57896
rect 1301 57838 1919 57840
rect 1301 57835 1367 57838
rect 1853 57835 1919 57838
rect 0 57762 800 57792
rect 2773 57762 2839 57765
rect 0 57760 2839 57762
rect 0 57704 2778 57760
rect 2834 57704 2839 57760
rect 0 57702 2839 57704
rect 0 57672 800 57702
rect 2773 57699 2839 57702
rect 4207 57696 4527 57697
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 4207 57631 4527 57632
rect 7471 57696 7791 57697
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 57631 7791 57632
rect 3182 57564 3188 57628
rect 3252 57626 3258 57628
rect 3693 57626 3759 57629
rect 3252 57624 3759 57626
rect 3252 57568 3698 57624
rect 3754 57568 3759 57624
rect 3252 57566 3759 57568
rect 3252 57564 3258 57566
rect 3693 57563 3759 57566
rect 1117 57490 1183 57493
rect 3233 57490 3299 57493
rect 1117 57488 3299 57490
rect 1117 57432 1122 57488
rect 1178 57432 3238 57488
rect 3294 57432 3299 57488
rect 1117 57430 3299 57432
rect 1117 57427 1183 57430
rect 3233 57427 3299 57430
rect 10133 57490 10199 57493
rect 11200 57490 12000 57520
rect 10133 57488 12000 57490
rect 10133 57432 10138 57488
rect 10194 57432 12000 57488
rect 10133 57430 12000 57432
rect 10133 57427 10199 57430
rect 11200 57400 12000 57430
rect 0 57354 800 57384
rect 1393 57354 1459 57357
rect 0 57352 1459 57354
rect 0 57296 1398 57352
rect 1454 57296 1459 57352
rect 0 57294 1459 57296
rect 0 57264 800 57294
rect 1393 57291 1459 57294
rect 2262 57292 2268 57356
rect 2332 57354 2338 57356
rect 2865 57354 2931 57357
rect 2332 57352 2931 57354
rect 2332 57296 2870 57352
rect 2926 57296 2931 57352
rect 2332 57294 2931 57296
rect 2332 57292 2338 57294
rect 2865 57291 2931 57294
rect 2576 57152 2896 57153
rect 2576 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2576 57087 2896 57088
rect 5839 57152 6159 57153
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 57087 6159 57088
rect 9103 57152 9423 57153
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 57087 9423 57088
rect 0 56946 800 56976
rect 1393 56946 1459 56949
rect 0 56944 1459 56946
rect 0 56888 1398 56944
rect 1454 56888 1459 56944
rect 0 56886 1459 56888
rect 0 56856 800 56886
rect 1393 56883 1459 56886
rect 10133 56674 10199 56677
rect 11200 56674 12000 56704
rect 10133 56672 12000 56674
rect 10133 56616 10138 56672
rect 10194 56616 12000 56672
rect 10133 56614 12000 56616
rect 10133 56611 10199 56614
rect 4207 56608 4527 56609
rect 0 56538 800 56568
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 4207 56543 4527 56544
rect 7471 56608 7791 56609
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 11200 56584 12000 56614
rect 7471 56543 7791 56544
rect 1485 56538 1551 56541
rect 0 56536 1551 56538
rect 0 56480 1490 56536
rect 1546 56480 1551 56536
rect 0 56478 1551 56480
rect 0 56448 800 56478
rect 1485 56475 1551 56478
rect 3141 56266 3207 56269
rect 3366 56266 3372 56268
rect 3141 56264 3372 56266
rect 3141 56208 3146 56264
rect 3202 56208 3372 56264
rect 3141 56206 3372 56208
rect 3141 56203 3207 56206
rect 3366 56204 3372 56206
rect 3436 56204 3442 56268
rect 2576 56064 2896 56065
rect 0 55994 800 56024
rect 2576 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2576 55999 2896 56000
rect 5839 56064 6159 56065
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 55999 6159 56000
rect 9103 56064 9423 56065
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 55999 9423 56000
rect 0 55934 1410 55994
rect 0 55904 800 55934
rect 1350 55858 1410 55934
rect 3141 55858 3207 55861
rect 1350 55856 3207 55858
rect 1350 55800 3146 55856
rect 3202 55800 3207 55856
rect 1350 55798 3207 55800
rect 3141 55795 3207 55798
rect 10133 55858 10199 55861
rect 11200 55858 12000 55888
rect 10133 55856 12000 55858
rect 10133 55800 10138 55856
rect 10194 55800 12000 55856
rect 10133 55798 12000 55800
rect 10133 55795 10199 55798
rect 11200 55768 12000 55798
rect 0 55586 800 55616
rect 3969 55586 4035 55589
rect 0 55584 4035 55586
rect 0 55528 3974 55584
rect 4030 55528 4035 55584
rect 0 55526 4035 55528
rect 0 55496 800 55526
rect 3969 55523 4035 55526
rect 4207 55520 4527 55521
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 55455 4527 55456
rect 7471 55520 7791 55521
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 55455 7791 55456
rect 3141 55452 3207 55453
rect 3141 55450 3188 55452
rect 3096 55448 3188 55450
rect 3096 55392 3146 55448
rect 3096 55390 3188 55392
rect 3141 55388 3188 55390
rect 3252 55388 3258 55452
rect 3141 55387 3207 55388
rect 0 55178 800 55208
rect 2773 55178 2839 55181
rect 0 55176 2839 55178
rect 0 55120 2778 55176
rect 2834 55120 2839 55176
rect 0 55118 2839 55120
rect 0 55088 800 55118
rect 2773 55115 2839 55118
rect 10133 55178 10199 55181
rect 11200 55178 12000 55208
rect 10133 55176 12000 55178
rect 10133 55120 10138 55176
rect 10194 55120 12000 55176
rect 10133 55118 12000 55120
rect 10133 55115 10199 55118
rect 11200 55088 12000 55118
rect 2576 54976 2896 54977
rect 2576 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2576 54911 2896 54912
rect 5839 54976 6159 54977
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 54911 6159 54912
rect 9103 54976 9423 54977
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 54911 9423 54912
rect 0 54770 800 54800
rect 1485 54770 1551 54773
rect 0 54768 1551 54770
rect 0 54712 1490 54768
rect 1546 54712 1551 54768
rect 0 54710 1551 54712
rect 0 54680 800 54710
rect 1485 54707 1551 54710
rect 1894 54572 1900 54636
rect 1964 54634 1970 54636
rect 2221 54634 2287 54637
rect 1964 54632 2287 54634
rect 1964 54576 2226 54632
rect 2282 54576 2287 54632
rect 1964 54574 2287 54576
rect 1964 54572 1970 54574
rect 2221 54571 2287 54574
rect 4207 54432 4527 54433
rect 0 54362 800 54392
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 54367 4527 54368
rect 7471 54432 7791 54433
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 54367 7791 54368
rect 2221 54362 2287 54365
rect 0 54360 2287 54362
rect 0 54304 2226 54360
rect 2282 54304 2287 54360
rect 0 54302 2287 54304
rect 0 54272 800 54302
rect 2221 54299 2287 54302
rect 10133 54362 10199 54365
rect 11200 54362 12000 54392
rect 10133 54360 12000 54362
rect 10133 54304 10138 54360
rect 10194 54304 12000 54360
rect 10133 54302 12000 54304
rect 10133 54299 10199 54302
rect 11200 54272 12000 54302
rect 0 53954 800 53984
rect 1485 53954 1551 53957
rect 0 53952 1551 53954
rect 0 53896 1490 53952
rect 1546 53896 1551 53952
rect 0 53894 1551 53896
rect 0 53864 800 53894
rect 1485 53891 1551 53894
rect 2576 53888 2896 53889
rect 2576 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2576 53823 2896 53824
rect 5839 53888 6159 53889
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 53823 6159 53824
rect 9103 53888 9423 53889
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 53823 9423 53824
rect 10041 53682 10107 53685
rect 11200 53682 12000 53712
rect 10041 53680 12000 53682
rect 10041 53624 10046 53680
rect 10102 53624 12000 53680
rect 10041 53622 12000 53624
rect 10041 53619 10107 53622
rect 11200 53592 12000 53622
rect 0 53546 800 53576
rect 2773 53546 2839 53549
rect 0 53544 2839 53546
rect 0 53488 2778 53544
rect 2834 53488 2839 53544
rect 0 53486 2839 53488
rect 0 53456 800 53486
rect 2773 53483 2839 53486
rect 4207 53344 4527 53345
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 53279 4527 53280
rect 7471 53344 7791 53345
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 53279 7791 53280
rect 0 53002 800 53032
rect 3049 53002 3115 53005
rect 0 53000 3115 53002
rect 0 52944 3054 53000
rect 3110 52944 3115 53000
rect 0 52942 3115 52944
rect 0 52912 800 52942
rect 3049 52939 3115 52942
rect 10041 52866 10107 52869
rect 11200 52866 12000 52896
rect 10041 52864 12000 52866
rect 10041 52808 10046 52864
rect 10102 52808 12000 52864
rect 10041 52806 12000 52808
rect 10041 52803 10107 52806
rect 2576 52800 2896 52801
rect 2576 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2576 52735 2896 52736
rect 5839 52800 6159 52801
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 52735 6159 52736
rect 9103 52800 9423 52801
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 11200 52776 12000 52806
rect 9103 52735 9423 52736
rect 0 52594 800 52624
rect 2221 52594 2287 52597
rect 0 52592 2287 52594
rect 0 52536 2226 52592
rect 2282 52536 2287 52592
rect 0 52534 2287 52536
rect 0 52504 800 52534
rect 2221 52531 2287 52534
rect 4207 52256 4527 52257
rect 0 52186 800 52216
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 4207 52191 4527 52192
rect 7471 52256 7791 52257
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 52191 7791 52192
rect 1393 52186 1459 52189
rect 0 52184 1459 52186
rect 0 52128 1398 52184
rect 1454 52128 1459 52184
rect 0 52126 1459 52128
rect 0 52096 800 52126
rect 1393 52123 1459 52126
rect 10041 52050 10107 52053
rect 11200 52050 12000 52080
rect 10041 52048 12000 52050
rect 10041 51992 10046 52048
rect 10102 51992 12000 52048
rect 10041 51990 12000 51992
rect 10041 51987 10107 51990
rect 11200 51960 12000 51990
rect 0 51778 800 51808
rect 1485 51778 1551 51781
rect 0 51776 1551 51778
rect 0 51720 1490 51776
rect 1546 51720 1551 51776
rect 0 51718 1551 51720
rect 0 51688 800 51718
rect 1485 51715 1551 51718
rect 2576 51712 2896 51713
rect 2576 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2576 51647 2896 51648
rect 5839 51712 6159 51713
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 51647 6159 51648
rect 9103 51712 9423 51713
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 51647 9423 51648
rect 0 51370 800 51400
rect 2221 51370 2287 51373
rect 0 51368 2287 51370
rect 0 51312 2226 51368
rect 2282 51312 2287 51368
rect 0 51310 2287 51312
rect 0 51280 800 51310
rect 2221 51307 2287 51310
rect 10041 51370 10107 51373
rect 11200 51370 12000 51400
rect 10041 51368 12000 51370
rect 10041 51312 10046 51368
rect 10102 51312 12000 51368
rect 10041 51310 12000 51312
rect 10041 51307 10107 51310
rect 11200 51280 12000 51310
rect 2129 51234 2195 51237
rect 1902 51232 2195 51234
rect 1902 51176 2134 51232
rect 2190 51176 2195 51232
rect 1902 51174 2195 51176
rect 1301 51090 1367 51093
rect 1301 51088 1410 51090
rect 1301 51032 1306 51088
rect 1362 51032 1410 51088
rect 1301 51027 1410 51032
rect 0 50962 800 50992
rect 1350 50962 1410 51027
rect 0 50902 1410 50962
rect 0 50872 800 50902
rect 1902 50826 1962 51174
rect 2129 51171 2195 51174
rect 3325 51234 3391 51237
rect 3918 51234 3924 51236
rect 3325 51232 3924 51234
rect 3325 51176 3330 51232
rect 3386 51176 3924 51232
rect 3325 51174 3924 51176
rect 3325 51171 3391 51174
rect 3918 51172 3924 51174
rect 3988 51172 3994 51236
rect 4207 51168 4527 51169
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 51103 4527 51104
rect 7471 51168 7791 51169
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 7471 51103 7791 51104
rect 2078 51036 2084 51100
rect 2148 51098 2154 51100
rect 2497 51098 2563 51101
rect 3693 51100 3759 51101
rect 3693 51098 3740 51100
rect 2148 51096 2563 51098
rect 2148 51040 2502 51096
rect 2558 51040 2563 51096
rect 2148 51038 2563 51040
rect 3648 51096 3740 51098
rect 3648 51040 3698 51096
rect 3648 51038 3740 51040
rect 2148 51036 2154 51038
rect 2497 51035 2563 51038
rect 3693 51036 3740 51038
rect 3804 51036 3810 51100
rect 3693 51035 3759 51036
rect 2221 50962 2287 50965
rect 2773 50962 2839 50965
rect 2221 50960 2839 50962
rect 2221 50904 2226 50960
rect 2282 50904 2778 50960
rect 2834 50904 2839 50960
rect 2221 50902 2839 50904
rect 2221 50899 2287 50902
rect 2773 50899 2839 50902
rect 3049 50962 3115 50965
rect 6310 50962 6316 50964
rect 3049 50960 6316 50962
rect 3049 50904 3054 50960
rect 3110 50904 6316 50960
rect 3049 50902 6316 50904
rect 3049 50899 3115 50902
rect 6310 50900 6316 50902
rect 6380 50900 6386 50964
rect 2129 50826 2195 50829
rect 1902 50824 2195 50826
rect 1902 50768 2134 50824
rect 2190 50768 2195 50824
rect 1902 50766 2195 50768
rect 2129 50763 2195 50766
rect 2262 50764 2268 50828
rect 2332 50826 2338 50828
rect 2497 50826 2563 50829
rect 2332 50824 2563 50826
rect 2332 50768 2502 50824
rect 2558 50768 2563 50824
rect 2332 50766 2563 50768
rect 2332 50764 2338 50766
rect 2497 50763 2563 50766
rect 2865 50826 2931 50829
rect 3325 50828 3391 50829
rect 2998 50826 3004 50828
rect 2865 50824 3004 50826
rect 2865 50768 2870 50824
rect 2926 50768 3004 50824
rect 2865 50766 3004 50768
rect 2865 50763 2931 50766
rect 2998 50764 3004 50766
rect 3068 50764 3074 50828
rect 3325 50824 3372 50828
rect 3436 50826 3442 50828
rect 3325 50768 3330 50824
rect 3325 50764 3372 50768
rect 3436 50766 3482 50826
rect 3436 50764 3442 50766
rect 3325 50763 3391 50764
rect 1894 50628 1900 50692
rect 1964 50690 1970 50692
rect 2037 50690 2103 50693
rect 1964 50688 2103 50690
rect 1964 50632 2042 50688
rect 2098 50632 2103 50688
rect 1964 50630 2103 50632
rect 1964 50628 1970 50630
rect 2037 50627 2103 50630
rect 2576 50624 2896 50625
rect 2576 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2576 50559 2896 50560
rect 5839 50624 6159 50625
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 5839 50559 6159 50560
rect 9103 50624 9423 50625
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 50559 9423 50560
rect 1301 50554 1367 50557
rect 798 50552 1367 50554
rect 798 50496 1306 50552
rect 1362 50496 1367 50552
rect 798 50494 1367 50496
rect 798 50448 858 50494
rect 1301 50491 1367 50494
rect 3182 50492 3188 50556
rect 3252 50554 3258 50556
rect 3785 50554 3851 50557
rect 3252 50552 3851 50554
rect 3252 50496 3790 50552
rect 3846 50496 3851 50552
rect 3252 50494 3851 50496
rect 3252 50492 3258 50494
rect 3785 50491 3851 50494
rect 10041 50554 10107 50557
rect 11200 50554 12000 50584
rect 10041 50552 12000 50554
rect 10041 50496 10046 50552
rect 10102 50496 12000 50552
rect 10041 50494 12000 50496
rect 10041 50491 10107 50494
rect 11200 50464 12000 50494
rect 0 50358 858 50448
rect 0 50328 800 50358
rect 4207 50080 4527 50081
rect 0 50010 800 50040
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 4207 50015 4527 50016
rect 7471 50080 7791 50081
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 7471 50015 7791 50016
rect 1485 50010 1551 50013
rect 0 50008 1551 50010
rect 0 49952 1490 50008
rect 1546 49952 1551 50008
rect 0 49950 1551 49952
rect 0 49920 800 49950
rect 1485 49947 1551 49950
rect 3918 49812 3924 49876
rect 3988 49874 3994 49876
rect 4153 49874 4219 49877
rect 3988 49872 4219 49874
rect 3988 49816 4158 49872
rect 4214 49816 4219 49872
rect 3988 49814 4219 49816
rect 3988 49812 3994 49814
rect 4153 49811 4219 49814
rect 10041 49874 10107 49877
rect 11200 49874 12000 49904
rect 10041 49872 12000 49874
rect 10041 49816 10046 49872
rect 10102 49816 12000 49872
rect 10041 49814 12000 49816
rect 10041 49811 10107 49814
rect 11200 49784 12000 49814
rect 2405 49738 2471 49741
rect 6494 49738 6500 49740
rect 2405 49736 6500 49738
rect 2405 49680 2410 49736
rect 2466 49680 6500 49736
rect 2405 49678 6500 49680
rect 2405 49675 2471 49678
rect 6494 49676 6500 49678
rect 6564 49676 6570 49740
rect 0 49602 800 49632
rect 2405 49602 2471 49605
rect 0 49600 2471 49602
rect 0 49544 2410 49600
rect 2466 49544 2471 49600
rect 0 49542 2471 49544
rect 0 49512 800 49542
rect 2405 49539 2471 49542
rect 3734 49540 3740 49604
rect 3804 49602 3810 49604
rect 3877 49602 3943 49605
rect 3804 49600 3943 49602
rect 3804 49544 3882 49600
rect 3938 49544 3943 49600
rect 3804 49542 3943 49544
rect 3804 49540 3810 49542
rect 3877 49539 3943 49542
rect 4654 49540 4660 49604
rect 4724 49602 4730 49604
rect 4797 49602 4863 49605
rect 4724 49600 4863 49602
rect 4724 49544 4802 49600
rect 4858 49544 4863 49600
rect 4724 49542 4863 49544
rect 4724 49540 4730 49542
rect 4797 49539 4863 49542
rect 2576 49536 2896 49537
rect 2576 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2576 49471 2896 49472
rect 5839 49536 6159 49537
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5839 49471 6159 49472
rect 9103 49536 9423 49537
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 49471 9423 49472
rect 0 49194 800 49224
rect 2221 49194 2287 49197
rect 0 49192 2287 49194
rect 0 49136 2226 49192
rect 2282 49136 2287 49192
rect 0 49134 2287 49136
rect 0 49104 800 49134
rect 2221 49131 2287 49134
rect 3877 49194 3943 49197
rect 6545 49194 6611 49197
rect 3877 49192 6611 49194
rect 3877 49136 3882 49192
rect 3938 49136 6550 49192
rect 6606 49136 6611 49192
rect 3877 49134 6611 49136
rect 3877 49131 3943 49134
rect 6545 49131 6611 49134
rect 1945 49058 2011 49061
rect 2078 49058 2084 49060
rect 1945 49056 2084 49058
rect 1945 49000 1950 49056
rect 2006 49000 2084 49056
rect 1945 48998 2084 49000
rect 1945 48995 2011 48998
rect 2078 48996 2084 48998
rect 2148 48996 2154 49060
rect 5390 48996 5396 49060
rect 5460 49058 5466 49060
rect 5625 49058 5691 49061
rect 5460 49056 5691 49058
rect 5460 49000 5630 49056
rect 5686 49000 5691 49056
rect 5460 48998 5691 49000
rect 5460 48996 5466 48998
rect 5625 48995 5691 48998
rect 10041 49058 10107 49061
rect 11200 49058 12000 49088
rect 10041 49056 12000 49058
rect 10041 49000 10046 49056
rect 10102 49000 12000 49056
rect 10041 48998 12000 49000
rect 10041 48995 10107 48998
rect 4207 48992 4527 48993
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 48927 4527 48928
rect 7471 48992 7791 48993
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 11200 48968 12000 48998
rect 7471 48927 7791 48928
rect 5533 48924 5599 48925
rect 5533 48920 5580 48924
rect 5644 48922 5650 48924
rect 5533 48864 5538 48920
rect 5533 48860 5580 48864
rect 5644 48862 5690 48922
rect 5644 48860 5650 48862
rect 5533 48859 5599 48860
rect 0 48786 800 48816
rect 2773 48786 2839 48789
rect 0 48784 2839 48786
rect 0 48728 2778 48784
rect 2834 48728 2839 48784
rect 0 48726 2839 48728
rect 0 48696 800 48726
rect 2773 48723 2839 48726
rect 2221 48650 2287 48653
rect 6821 48650 6887 48653
rect 2221 48648 6887 48650
rect 2221 48592 2226 48648
rect 2282 48592 6826 48648
rect 6882 48592 6887 48648
rect 2221 48590 6887 48592
rect 2221 48587 2287 48590
rect 6821 48587 6887 48590
rect 5390 48452 5396 48516
rect 5460 48514 5466 48516
rect 5625 48514 5691 48517
rect 5460 48512 5691 48514
rect 5460 48456 5630 48512
rect 5686 48456 5691 48512
rect 5460 48454 5691 48456
rect 5460 48452 5466 48454
rect 5625 48451 5691 48454
rect 2576 48448 2896 48449
rect 0 48378 800 48408
rect 2576 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2576 48383 2896 48384
rect 5839 48448 6159 48449
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5839 48383 6159 48384
rect 9103 48448 9423 48449
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 48383 9423 48384
rect 1485 48378 1551 48381
rect 0 48376 1551 48378
rect 0 48320 1490 48376
rect 1546 48320 1551 48376
rect 5574 48347 5580 48380
rect 5533 48344 5580 48347
rect 0 48318 1551 48320
rect 0 48288 800 48318
rect 1485 48315 1551 48318
rect 5522 48342 5580 48344
rect 5522 48286 5538 48342
rect 5644 48316 5650 48380
rect 5594 48286 5642 48316
rect 5522 48284 5642 48286
rect 5533 48281 5599 48284
rect 2262 48180 2268 48244
rect 2332 48242 2338 48244
rect 2681 48242 2747 48245
rect 2332 48240 2747 48242
rect 2332 48184 2686 48240
rect 2742 48184 2747 48240
rect 2332 48182 2747 48184
rect 2332 48180 2338 48182
rect 2681 48179 2747 48182
rect 10041 48242 10107 48245
rect 11200 48242 12000 48272
rect 10041 48240 12000 48242
rect 10041 48184 10046 48240
rect 10102 48184 12000 48240
rect 10041 48182 12000 48184
rect 10041 48179 10107 48182
rect 11200 48152 12000 48182
rect 4207 47904 4527 47905
rect 0 47834 800 47864
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 47839 4527 47840
rect 7471 47904 7791 47905
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 47839 7791 47840
rect 1485 47834 1551 47837
rect 0 47832 1551 47834
rect 0 47776 1490 47832
rect 1546 47776 1551 47832
rect 0 47774 1551 47776
rect 0 47744 800 47774
rect 1485 47771 1551 47774
rect 4838 47772 4844 47836
rect 4908 47834 4914 47836
rect 6177 47834 6243 47837
rect 4908 47832 6243 47834
rect 4908 47776 6182 47832
rect 6238 47776 6243 47832
rect 4908 47774 6243 47776
rect 4908 47772 4914 47774
rect 6177 47771 6243 47774
rect 10041 47562 10107 47565
rect 11200 47562 12000 47592
rect 10041 47560 12000 47562
rect 10041 47504 10046 47560
rect 10102 47504 12000 47560
rect 10041 47502 12000 47504
rect 10041 47499 10107 47502
rect 11200 47472 12000 47502
rect 0 47426 800 47456
rect 2221 47426 2287 47429
rect 0 47424 2287 47426
rect 0 47368 2226 47424
rect 2282 47368 2287 47424
rect 0 47366 2287 47368
rect 0 47336 800 47366
rect 2221 47363 2287 47366
rect 2576 47360 2896 47361
rect 2576 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2576 47295 2896 47296
rect 5839 47360 6159 47361
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 47295 6159 47296
rect 9103 47360 9423 47361
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 47295 9423 47296
rect 0 47018 800 47048
rect 1485 47018 1551 47021
rect 0 47016 1551 47018
rect 0 46960 1490 47016
rect 1546 46960 1551 47016
rect 0 46958 1551 46960
rect 0 46928 800 46958
rect 1485 46955 1551 46958
rect 4207 46816 4527 46817
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 4207 46751 4527 46752
rect 7471 46816 7791 46817
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 46751 7791 46752
rect 3049 46746 3115 46749
rect 3182 46746 3188 46748
rect 3049 46744 3188 46746
rect 3049 46688 3054 46744
rect 3110 46688 3188 46744
rect 3049 46686 3188 46688
rect 3049 46683 3115 46686
rect 3182 46684 3188 46686
rect 3252 46684 3258 46748
rect 10041 46746 10107 46749
rect 11200 46746 12000 46776
rect 10041 46744 12000 46746
rect 10041 46688 10046 46744
rect 10102 46688 12000 46744
rect 10041 46686 12000 46688
rect 10041 46683 10107 46686
rect 11200 46656 12000 46686
rect 0 46610 800 46640
rect 1485 46610 1551 46613
rect 0 46608 1551 46610
rect 0 46552 1490 46608
rect 1546 46552 1551 46608
rect 0 46550 1551 46552
rect 0 46520 800 46550
rect 1485 46547 1551 46550
rect 2313 46474 2379 46477
rect 3918 46474 3924 46476
rect 2313 46472 3924 46474
rect 2313 46416 2318 46472
rect 2374 46416 3924 46472
rect 2313 46414 3924 46416
rect 2313 46411 2379 46414
rect 3918 46412 3924 46414
rect 3988 46412 3994 46476
rect 6453 46474 6519 46477
rect 7005 46474 7071 46477
rect 6453 46472 6746 46474
rect 6453 46416 6458 46472
rect 6514 46416 6746 46472
rect 6453 46414 6746 46416
rect 6453 46411 6519 46414
rect 2576 46272 2896 46273
rect 0 46202 800 46232
rect 2576 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2576 46207 2896 46208
rect 5839 46272 6159 46273
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5839 46207 6159 46208
rect 1485 46202 1551 46205
rect 0 46200 1551 46202
rect 0 46144 1490 46200
rect 1546 46144 1551 46200
rect 0 46142 1551 46144
rect 0 46112 800 46142
rect 1485 46139 1551 46142
rect 4889 46202 4955 46205
rect 5022 46202 5028 46204
rect 4889 46200 5028 46202
rect 4889 46144 4894 46200
rect 4950 46144 5028 46200
rect 4889 46142 5028 46144
rect 4889 46139 4955 46142
rect 5022 46140 5028 46142
rect 5092 46140 5098 46204
rect 6686 46069 6746 46414
rect 6870 46472 7071 46474
rect 6870 46416 7010 46472
rect 7066 46416 7071 46472
rect 6870 46414 7071 46416
rect 2129 46066 2195 46069
rect 2998 46066 3004 46068
rect 2129 46064 3004 46066
rect 2129 46008 2134 46064
rect 2190 46008 3004 46064
rect 2129 46006 3004 46008
rect 2129 46003 2195 46006
rect 2998 46004 3004 46006
rect 3068 46004 3074 46068
rect 6686 46064 6795 46069
rect 6686 46008 6734 46064
rect 6790 46008 6795 46064
rect 6686 46006 6795 46008
rect 6729 46003 6795 46006
rect 5717 45930 5783 45933
rect 6870 45930 6930 46414
rect 7005 46411 7071 46414
rect 7925 46474 7991 46477
rect 7925 46472 8034 46474
rect 7925 46416 7930 46472
rect 7986 46416 8034 46472
rect 7925 46411 8034 46416
rect 7974 46066 8034 46411
rect 9103 46272 9423 46273
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 46207 9423 46208
rect 8109 46066 8175 46069
rect 7974 46064 8175 46066
rect 7974 46008 8114 46064
rect 8170 46008 8175 46064
rect 7974 46006 8175 46008
rect 8109 46003 8175 46006
rect 10041 46066 10107 46069
rect 11200 46066 12000 46096
rect 10041 46064 12000 46066
rect 10041 46008 10046 46064
rect 10102 46008 12000 46064
rect 10041 46006 12000 46008
rect 10041 46003 10107 46006
rect 11200 45976 12000 46006
rect 5717 45928 6930 45930
rect 5717 45872 5722 45928
rect 5778 45872 6930 45928
rect 5717 45870 6930 45872
rect 5717 45867 5783 45870
rect 0 45794 800 45824
rect 2957 45794 3023 45797
rect 0 45792 3023 45794
rect 0 45736 2962 45792
rect 3018 45736 3023 45792
rect 0 45734 3023 45736
rect 0 45704 800 45734
rect 2957 45731 3023 45734
rect 4207 45728 4527 45729
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 45663 4527 45664
rect 7471 45728 7791 45729
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 45663 7791 45664
rect 2405 45658 2471 45661
rect 3417 45658 3483 45661
rect 2405 45656 3483 45658
rect 2405 45600 2410 45656
rect 2466 45600 3422 45656
rect 3478 45600 3483 45656
rect 2405 45598 3483 45600
rect 2405 45595 2471 45598
rect 3417 45595 3483 45598
rect 0 45250 800 45280
rect 1485 45250 1551 45253
rect 0 45248 1551 45250
rect 0 45192 1490 45248
rect 1546 45192 1551 45248
rect 0 45190 1551 45192
rect 0 45160 800 45190
rect 1485 45187 1551 45190
rect 10041 45250 10107 45253
rect 11200 45250 12000 45280
rect 10041 45248 12000 45250
rect 10041 45192 10046 45248
rect 10102 45192 12000 45248
rect 10041 45190 12000 45192
rect 10041 45187 10107 45190
rect 2576 45184 2896 45185
rect 2576 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2576 45119 2896 45120
rect 5839 45184 6159 45185
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 45119 6159 45120
rect 9103 45184 9423 45185
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 11200 45160 12000 45190
rect 9103 45119 9423 45120
rect 2037 45116 2103 45117
rect 2037 45112 2084 45116
rect 2148 45114 2154 45116
rect 2037 45056 2042 45112
rect 2037 45052 2084 45056
rect 2148 45054 2194 45114
rect 2148 45052 2154 45054
rect 2998 45052 3004 45116
rect 3068 45114 3074 45116
rect 4981 45114 5047 45117
rect 3068 45112 5047 45114
rect 3068 45056 4986 45112
rect 5042 45056 5047 45112
rect 3068 45054 5047 45056
rect 3068 45052 3074 45054
rect 2037 45051 2103 45052
rect 4981 45051 5047 45054
rect 3785 44978 3851 44981
rect 3742 44976 3851 44978
rect 3742 44920 3790 44976
rect 3846 44920 3851 44976
rect 3742 44915 3851 44920
rect 0 44842 800 44872
rect 2405 44842 2471 44845
rect 0 44840 2471 44842
rect 0 44784 2410 44840
rect 2466 44784 2471 44840
rect 0 44782 2471 44784
rect 0 44752 800 44782
rect 2405 44779 2471 44782
rect 0 44434 800 44464
rect 1577 44434 1643 44437
rect 0 44432 1643 44434
rect 0 44376 1582 44432
rect 1638 44376 1643 44432
rect 0 44374 1643 44376
rect 0 44344 800 44374
rect 1577 44371 1643 44374
rect 3601 44434 3667 44437
rect 3742 44434 3802 44915
rect 4207 44640 4527 44641
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 44575 4527 44576
rect 7471 44640 7791 44641
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 44575 7791 44576
rect 3601 44432 3802 44434
rect 3601 44376 3606 44432
rect 3662 44376 3802 44432
rect 3601 44374 3802 44376
rect 10041 44434 10107 44437
rect 11200 44434 12000 44464
rect 10041 44432 12000 44434
rect 10041 44376 10046 44432
rect 10102 44376 12000 44432
rect 10041 44374 12000 44376
rect 3601 44371 3667 44374
rect 10041 44371 10107 44374
rect 11200 44344 12000 44374
rect 2576 44096 2896 44097
rect 0 44026 800 44056
rect 2576 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2576 44031 2896 44032
rect 5839 44096 6159 44097
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 44031 6159 44032
rect 9103 44096 9423 44097
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 44031 9423 44032
rect 2405 44026 2471 44029
rect 0 44024 2471 44026
rect 0 43968 2410 44024
rect 2466 43968 2471 44024
rect 0 43966 2471 43968
rect 0 43936 800 43966
rect 2405 43963 2471 43966
rect 10041 43754 10107 43757
rect 11200 43754 12000 43784
rect 10041 43752 12000 43754
rect 10041 43696 10046 43752
rect 10102 43696 12000 43752
rect 10041 43694 12000 43696
rect 10041 43691 10107 43694
rect 11200 43664 12000 43694
rect 0 43618 800 43648
rect 3049 43618 3115 43621
rect 0 43616 3115 43618
rect 0 43560 3054 43616
rect 3110 43560 3115 43616
rect 0 43558 3115 43560
rect 0 43528 800 43558
rect 3049 43555 3115 43558
rect 4207 43552 4527 43553
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 43487 4527 43488
rect 7471 43552 7791 43553
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 43487 7791 43488
rect 2313 43484 2379 43485
rect 2262 43482 2268 43484
rect 2222 43422 2268 43482
rect 2332 43480 2379 43484
rect 2374 43424 2379 43480
rect 2262 43420 2268 43422
rect 2332 43420 2379 43424
rect 2313 43419 2379 43420
rect 2865 43346 2931 43349
rect 3049 43346 3115 43349
rect 3182 43346 3188 43348
rect 2865 43344 3188 43346
rect 2865 43288 2870 43344
rect 2926 43288 3054 43344
rect 3110 43288 3188 43344
rect 2865 43286 3188 43288
rect 2865 43283 2931 43286
rect 3049 43283 3115 43286
rect 3182 43284 3188 43286
rect 3252 43284 3258 43348
rect 4521 43346 4587 43349
rect 4654 43346 4660 43348
rect 4521 43344 4660 43346
rect 4521 43288 4526 43344
rect 4582 43288 4660 43344
rect 4521 43286 4660 43288
rect 4521 43283 4587 43286
rect 4654 43284 4660 43286
rect 4724 43284 4730 43348
rect 0 43210 800 43240
rect 2221 43210 2287 43213
rect 0 43208 2287 43210
rect 0 43152 2226 43208
rect 2282 43152 2287 43208
rect 0 43150 2287 43152
rect 0 43120 800 43150
rect 2221 43147 2287 43150
rect 2576 43008 2896 43009
rect 2576 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2576 42943 2896 42944
rect 5839 43008 6159 43009
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5839 42943 6159 42944
rect 9103 43008 9423 43009
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 42943 9423 42944
rect 10041 42938 10107 42941
rect 11200 42938 12000 42968
rect 10041 42936 12000 42938
rect 10041 42880 10046 42936
rect 10102 42880 12000 42936
rect 10041 42878 12000 42880
rect 10041 42875 10107 42878
rect 11200 42848 12000 42878
rect 0 42666 800 42696
rect 2221 42666 2287 42669
rect 0 42664 2287 42666
rect 0 42608 2226 42664
rect 2282 42608 2287 42664
rect 0 42606 2287 42608
rect 0 42576 800 42606
rect 2221 42603 2287 42606
rect 4207 42464 4527 42465
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 42399 4527 42400
rect 7471 42464 7791 42465
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 42399 7791 42400
rect 0 42258 800 42288
rect 1485 42258 1551 42261
rect 0 42256 1551 42258
rect 0 42200 1490 42256
rect 1546 42200 1551 42256
rect 0 42198 1551 42200
rect 0 42168 800 42198
rect 1485 42195 1551 42198
rect 1853 42258 1919 42261
rect 4153 42258 4219 42261
rect 4838 42258 4844 42260
rect 1853 42256 1962 42258
rect 1853 42200 1858 42256
rect 1914 42200 1962 42256
rect 1853 42195 1962 42200
rect 4153 42256 4844 42258
rect 4153 42200 4158 42256
rect 4214 42200 4844 42256
rect 4153 42198 4844 42200
rect 4153 42195 4219 42198
rect 4838 42196 4844 42198
rect 4908 42196 4914 42260
rect 10041 42258 10107 42261
rect 11200 42258 12000 42288
rect 10041 42256 12000 42258
rect 10041 42200 10046 42256
rect 10102 42200 12000 42256
rect 10041 42198 12000 42200
rect 10041 42195 10107 42198
rect 0 41850 800 41880
rect 1902 41853 1962 42195
rect 11200 42168 12000 42198
rect 2037 42124 2103 42125
rect 2037 42120 2084 42124
rect 2148 42122 2154 42124
rect 2037 42064 2042 42120
rect 2037 42060 2084 42064
rect 2148 42062 2194 42122
rect 2148 42060 2154 42062
rect 2037 42059 2103 42060
rect 5073 41988 5139 41989
rect 5022 41986 5028 41988
rect 4982 41926 5028 41986
rect 5092 41984 5139 41988
rect 5134 41928 5139 41984
rect 5022 41924 5028 41926
rect 5092 41924 5139 41928
rect 5073 41923 5139 41924
rect 2576 41920 2896 41921
rect 2576 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2576 41855 2896 41856
rect 5839 41920 6159 41921
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5839 41855 6159 41856
rect 9103 41920 9423 41921
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 41855 9423 41856
rect 1393 41850 1459 41853
rect 0 41848 1459 41850
rect 0 41792 1398 41848
rect 1454 41792 1459 41848
rect 0 41790 1459 41792
rect 0 41760 800 41790
rect 1393 41787 1459 41790
rect 1853 41848 1962 41853
rect 1853 41792 1858 41848
rect 1914 41792 1962 41848
rect 1853 41790 1962 41792
rect 1853 41787 1919 41790
rect 4797 41714 4863 41717
rect 5390 41714 5396 41716
rect 4797 41712 5396 41714
rect 4797 41656 4802 41712
rect 4858 41656 5396 41712
rect 4797 41654 5396 41656
rect 4797 41651 4863 41654
rect 5390 41652 5396 41654
rect 5460 41652 5466 41716
rect 5206 41516 5212 41580
rect 5276 41578 5282 41580
rect 5349 41578 5415 41581
rect 5276 41576 5415 41578
rect 5276 41520 5354 41576
rect 5410 41520 5415 41576
rect 5276 41518 5415 41520
rect 5276 41516 5282 41518
rect 5349 41515 5415 41518
rect 6177 41578 6243 41581
rect 6310 41578 6316 41580
rect 6177 41576 6316 41578
rect 6177 41520 6182 41576
rect 6238 41520 6316 41576
rect 6177 41518 6316 41520
rect 6177 41515 6243 41518
rect 6310 41516 6316 41518
rect 6380 41516 6386 41580
rect 6729 41578 6795 41581
rect 6686 41576 6795 41578
rect 6686 41520 6734 41576
rect 6790 41520 6795 41576
rect 6686 41515 6795 41520
rect 0 41442 800 41472
rect 1485 41442 1551 41445
rect 0 41440 1551 41442
rect 0 41384 1490 41440
rect 1546 41384 1551 41440
rect 0 41382 1551 41384
rect 0 41352 800 41382
rect 1485 41379 1551 41382
rect 6453 41442 6519 41445
rect 6686 41442 6746 41515
rect 6453 41440 6746 41442
rect 6453 41384 6458 41440
rect 6514 41384 6746 41440
rect 6453 41382 6746 41384
rect 10041 41442 10107 41445
rect 11200 41442 12000 41472
rect 10041 41440 12000 41442
rect 10041 41384 10046 41440
rect 10102 41384 12000 41440
rect 10041 41382 12000 41384
rect 6453 41379 6519 41382
rect 10041 41379 10107 41382
rect 4207 41376 4527 41377
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 41311 4527 41312
rect 7471 41376 7791 41377
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 11200 41352 12000 41382
rect 7471 41311 7791 41312
rect 1761 41306 1827 41309
rect 2129 41306 2195 41309
rect 2313 41308 2379 41309
rect 1761 41304 2195 41306
rect 1761 41248 1766 41304
rect 1822 41248 2134 41304
rect 2190 41248 2195 41304
rect 1761 41246 2195 41248
rect 1761 41243 1827 41246
rect 2129 41243 2195 41246
rect 2262 41244 2268 41308
rect 2332 41306 2379 41308
rect 2332 41304 2424 41306
rect 2374 41248 2424 41304
rect 2332 41246 2424 41248
rect 2332 41244 2379 41246
rect 6494 41244 6500 41308
rect 6564 41306 6570 41308
rect 6729 41306 6795 41309
rect 6564 41304 6795 41306
rect 6564 41248 6734 41304
rect 6790 41248 6795 41304
rect 6564 41246 6795 41248
rect 6564 41244 6570 41246
rect 2313 41243 2379 41244
rect 6729 41243 6795 41246
rect 1158 41108 1164 41172
rect 1228 41170 1234 41172
rect 1669 41170 1735 41173
rect 1228 41168 1735 41170
rect 1228 41112 1674 41168
rect 1730 41112 1735 41168
rect 1228 41110 1735 41112
rect 1228 41108 1234 41110
rect 1669 41107 1735 41110
rect 0 41034 800 41064
rect 2313 41034 2379 41037
rect 0 41032 2379 41034
rect 0 40976 2318 41032
rect 2374 40976 2379 41032
rect 0 40974 2379 40976
rect 0 40944 800 40974
rect 2313 40971 2379 40974
rect 2576 40832 2896 40833
rect 2576 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2576 40767 2896 40768
rect 5839 40832 6159 40833
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 40767 6159 40768
rect 9103 40832 9423 40833
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 40767 9423 40768
rect 0 40626 800 40656
rect 1393 40626 1459 40629
rect 0 40624 1459 40626
rect 0 40568 1398 40624
rect 1454 40568 1459 40624
rect 0 40566 1459 40568
rect 0 40536 800 40566
rect 1393 40563 1459 40566
rect 10041 40626 10107 40629
rect 11200 40626 12000 40656
rect 10041 40624 12000 40626
rect 10041 40568 10046 40624
rect 10102 40568 12000 40624
rect 10041 40566 12000 40568
rect 10041 40563 10107 40566
rect 11200 40536 12000 40566
rect 4207 40288 4527 40289
rect 0 40218 800 40248
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 40223 4527 40224
rect 7471 40288 7791 40289
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 40223 7791 40224
rect 3049 40218 3115 40221
rect 0 40216 3115 40218
rect 0 40160 3054 40216
rect 3110 40160 3115 40216
rect 0 40158 3115 40160
rect 0 40128 800 40158
rect 3049 40155 3115 40158
rect 4061 40082 4127 40085
rect 3742 40080 4127 40082
rect 3742 40024 4066 40080
rect 4122 40024 4127 40080
rect 3742 40022 4127 40024
rect 3509 39946 3575 39949
rect 3742 39946 3802 40022
rect 4061 40019 4127 40022
rect 3509 39944 3802 39946
rect 3509 39888 3514 39944
rect 3570 39888 3802 39944
rect 3509 39886 3802 39888
rect 10041 39946 10107 39949
rect 11200 39946 12000 39976
rect 10041 39944 12000 39946
rect 10041 39888 10046 39944
rect 10102 39888 12000 39944
rect 10041 39886 12000 39888
rect 3509 39883 3575 39886
rect 10041 39883 10107 39886
rect 11200 39856 12000 39886
rect 5165 39812 5231 39813
rect 5165 39810 5212 39812
rect 5120 39808 5212 39810
rect 5120 39752 5170 39808
rect 5120 39750 5212 39752
rect 5165 39748 5212 39750
rect 5276 39748 5282 39812
rect 5165 39747 5231 39748
rect 2576 39744 2896 39745
rect 0 39674 800 39704
rect 2576 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2576 39679 2896 39680
rect 5839 39744 6159 39745
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5839 39679 6159 39680
rect 9103 39744 9423 39745
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 39679 9423 39680
rect 2313 39674 2379 39677
rect 0 39672 2379 39674
rect 0 39616 2318 39672
rect 2374 39616 2379 39672
rect 0 39614 2379 39616
rect 0 39584 800 39614
rect 2313 39611 2379 39614
rect 3877 39538 3943 39541
rect 4889 39538 4955 39541
rect 5390 39538 5396 39540
rect 3877 39536 3986 39538
rect 3877 39480 3882 39536
rect 3938 39480 3986 39536
rect 3877 39475 3986 39480
rect 4889 39536 5396 39538
rect 4889 39480 4894 39536
rect 4950 39480 5396 39536
rect 4889 39478 5396 39480
rect 4889 39475 4955 39478
rect 5390 39476 5396 39478
rect 5460 39476 5466 39540
rect 0 39266 800 39296
rect 1485 39266 1551 39269
rect 0 39264 1551 39266
rect 0 39208 1490 39264
rect 1546 39208 1551 39264
rect 0 39206 1551 39208
rect 0 39176 800 39206
rect 1485 39203 1551 39206
rect 3926 38994 3986 39475
rect 4207 39200 4527 39201
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 4207 39135 4527 39136
rect 7471 39200 7791 39201
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 39135 7791 39136
rect 10041 39130 10107 39133
rect 11200 39130 12000 39160
rect 10041 39128 12000 39130
rect 10041 39072 10046 39128
rect 10102 39072 12000 39128
rect 10041 39070 12000 39072
rect 10041 39067 10107 39070
rect 11200 39040 12000 39070
rect 4061 38994 4127 38997
rect 3926 38992 4127 38994
rect 3926 38936 4066 38992
rect 4122 38936 4127 38992
rect 3926 38934 4127 38936
rect 4061 38931 4127 38934
rect 0 38858 800 38888
rect 2957 38858 3023 38861
rect 0 38856 3023 38858
rect 0 38800 2962 38856
rect 3018 38800 3023 38856
rect 0 38798 3023 38800
rect 0 38768 800 38798
rect 2957 38795 3023 38798
rect 3918 38796 3924 38860
rect 3988 38858 3994 38860
rect 4337 38858 4403 38861
rect 3988 38856 4403 38858
rect 3988 38800 4342 38856
rect 4398 38800 4403 38856
rect 3988 38798 4403 38800
rect 3988 38796 3994 38798
rect 4337 38795 4403 38798
rect 2078 38660 2084 38724
rect 2148 38722 2154 38724
rect 2405 38722 2471 38725
rect 2148 38720 2471 38722
rect 2148 38664 2410 38720
rect 2466 38664 2471 38720
rect 2148 38662 2471 38664
rect 2148 38660 2154 38662
rect 2405 38659 2471 38662
rect 2957 38724 3023 38725
rect 2957 38720 3004 38724
rect 3068 38722 3074 38724
rect 2957 38664 2962 38720
rect 2957 38660 3004 38664
rect 3068 38662 3114 38722
rect 3068 38660 3074 38662
rect 2957 38659 3023 38660
rect 2576 38656 2896 38657
rect 2576 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2576 38591 2896 38592
rect 5839 38656 6159 38657
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 38591 6159 38592
rect 9103 38656 9423 38657
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 38591 9423 38592
rect 0 38450 800 38480
rect 2221 38450 2287 38453
rect 0 38448 2287 38450
rect 0 38392 2226 38448
rect 2282 38392 2287 38448
rect 0 38390 2287 38392
rect 0 38360 800 38390
rect 2221 38387 2287 38390
rect 10041 38450 10107 38453
rect 11200 38450 12000 38480
rect 10041 38448 12000 38450
rect 10041 38392 10046 38448
rect 10102 38392 12000 38448
rect 10041 38390 12000 38392
rect 10041 38387 10107 38390
rect 11200 38360 12000 38390
rect 4207 38112 4527 38113
rect 0 38042 800 38072
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 4207 38047 4527 38048
rect 7471 38112 7791 38113
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 38047 7791 38048
rect 1393 38042 1459 38045
rect 0 38040 1459 38042
rect 0 37984 1398 38040
rect 1454 37984 1459 38040
rect 0 37982 1459 37984
rect 0 37952 800 37982
rect 1393 37979 1459 37982
rect 0 37634 800 37664
rect 2313 37634 2379 37637
rect 0 37632 2379 37634
rect 0 37576 2318 37632
rect 2374 37576 2379 37632
rect 0 37574 2379 37576
rect 0 37544 800 37574
rect 2313 37571 2379 37574
rect 10041 37634 10107 37637
rect 11200 37634 12000 37664
rect 10041 37632 12000 37634
rect 10041 37576 10046 37632
rect 10102 37576 12000 37632
rect 10041 37574 12000 37576
rect 10041 37571 10107 37574
rect 2576 37568 2896 37569
rect 2576 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2576 37503 2896 37504
rect 5839 37568 6159 37569
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 37503 6159 37504
rect 9103 37568 9423 37569
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 11200 37544 12000 37574
rect 9103 37503 9423 37504
rect 3734 37300 3740 37364
rect 3804 37362 3810 37364
rect 3969 37362 4035 37365
rect 3804 37360 4035 37362
rect 3804 37304 3974 37360
rect 4030 37304 4035 37360
rect 3804 37302 4035 37304
rect 3804 37300 3810 37302
rect 3969 37299 4035 37302
rect 2957 37228 3023 37229
rect 2957 37226 3004 37228
rect 2912 37224 3004 37226
rect 2912 37168 2962 37224
rect 2912 37166 3004 37168
rect 2957 37164 3004 37166
rect 3068 37164 3074 37228
rect 2957 37163 3023 37164
rect 0 37090 800 37120
rect 1485 37090 1551 37093
rect 0 37088 1551 37090
rect 0 37032 1490 37088
rect 1546 37032 1551 37088
rect 0 37030 1551 37032
rect 0 37000 800 37030
rect 1485 37027 1551 37030
rect 4207 37024 4527 37025
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 36959 4527 36960
rect 7471 37024 7791 37025
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 36959 7791 36960
rect 3509 36954 3575 36957
rect 3877 36954 3943 36957
rect 3509 36952 3943 36954
rect 3509 36896 3514 36952
rect 3570 36896 3882 36952
rect 3938 36896 3943 36952
rect 3509 36894 3943 36896
rect 3509 36891 3575 36894
rect 3877 36891 3943 36894
rect 10041 36818 10107 36821
rect 11200 36818 12000 36848
rect 10041 36816 12000 36818
rect 10041 36760 10046 36816
rect 10102 36760 12000 36816
rect 10041 36758 12000 36760
rect 10041 36755 10107 36758
rect 11200 36728 12000 36758
rect 0 36682 800 36712
rect 3049 36682 3115 36685
rect 3509 36684 3575 36685
rect 3509 36682 3556 36684
rect 0 36680 3115 36682
rect 0 36624 3054 36680
rect 3110 36624 3115 36680
rect 0 36622 3115 36624
rect 3464 36680 3556 36682
rect 3464 36624 3514 36680
rect 3464 36622 3556 36624
rect 0 36592 800 36622
rect 3049 36619 3115 36622
rect 3509 36620 3556 36622
rect 3620 36620 3626 36684
rect 7925 36682 7991 36685
rect 7925 36680 8034 36682
rect 7925 36624 7930 36680
rect 7986 36624 8034 36680
rect 3509 36619 3575 36620
rect 7925 36619 8034 36624
rect 2576 36480 2896 36481
rect 2576 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2576 36415 2896 36416
rect 5839 36480 6159 36481
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 36415 6159 36416
rect 5073 36410 5139 36413
rect 5257 36410 5323 36413
rect 5073 36408 5323 36410
rect 5073 36352 5078 36408
rect 5134 36352 5262 36408
rect 5318 36352 5323 36408
rect 5073 36350 5323 36352
rect 7974 36410 8034 36619
rect 9103 36480 9423 36481
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 36415 9423 36416
rect 8109 36410 8175 36413
rect 7974 36408 8175 36410
rect 7974 36352 8114 36408
rect 8170 36352 8175 36408
rect 7974 36350 8175 36352
rect 5073 36347 5139 36350
rect 5257 36347 5323 36350
rect 8109 36347 8175 36350
rect 0 36274 800 36304
rect 2221 36274 2287 36277
rect 0 36272 2287 36274
rect 0 36216 2226 36272
rect 2282 36216 2287 36272
rect 0 36214 2287 36216
rect 0 36184 800 36214
rect 2221 36211 2287 36214
rect 1485 36140 1551 36141
rect 1485 36138 1532 36140
rect 1440 36136 1532 36138
rect 1440 36080 1490 36136
rect 1440 36078 1532 36080
rect 1485 36076 1532 36078
rect 1596 36076 1602 36140
rect 10041 36138 10107 36141
rect 11200 36138 12000 36168
rect 10041 36136 12000 36138
rect 10041 36080 10046 36136
rect 10102 36080 12000 36136
rect 10041 36078 12000 36080
rect 1485 36075 1551 36076
rect 10041 36075 10107 36078
rect 11200 36048 12000 36078
rect 4207 35936 4527 35937
rect 0 35866 800 35896
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 4207 35871 4527 35872
rect 7471 35936 7791 35937
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 35871 7791 35872
rect 1393 35866 1459 35869
rect 0 35864 1459 35866
rect 0 35808 1398 35864
rect 1454 35808 1459 35864
rect 0 35806 1459 35808
rect 0 35776 800 35806
rect 1393 35803 1459 35806
rect 2405 35864 2471 35869
rect 2405 35808 2410 35864
rect 2466 35808 2471 35864
rect 2405 35803 2471 35808
rect 1393 35730 1459 35733
rect 2408 35730 2468 35803
rect 1393 35728 2468 35730
rect 1393 35672 1398 35728
rect 1454 35672 2468 35728
rect 1393 35670 2468 35672
rect 1393 35667 1459 35670
rect 4981 35594 5047 35597
rect 4981 35592 5274 35594
rect 4981 35536 4986 35592
rect 5042 35536 5274 35592
rect 4981 35534 5274 35536
rect 4981 35531 5047 35534
rect 0 35458 800 35488
rect 1485 35458 1551 35461
rect 0 35456 1551 35458
rect 0 35400 1490 35456
rect 1546 35400 1551 35456
rect 0 35398 1551 35400
rect 0 35368 800 35398
rect 1485 35395 1551 35398
rect 3693 35460 3759 35461
rect 3693 35456 3740 35460
rect 3804 35458 3810 35460
rect 3693 35400 3698 35456
rect 3693 35396 3740 35400
rect 3804 35398 3850 35458
rect 3804 35396 3810 35398
rect 3693 35395 3759 35396
rect 2576 35392 2896 35393
rect 2576 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2576 35327 2896 35328
rect 5214 35189 5274 35534
rect 5839 35392 6159 35393
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 35327 6159 35328
rect 9103 35392 9423 35393
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 35327 9423 35328
rect 10041 35322 10107 35325
rect 11200 35322 12000 35352
rect 10041 35320 12000 35322
rect 10041 35264 10046 35320
rect 10102 35264 12000 35320
rect 10041 35262 12000 35264
rect 10041 35259 10107 35262
rect 11200 35232 12000 35262
rect 5214 35184 5323 35189
rect 5214 35128 5262 35184
rect 5318 35128 5323 35184
rect 5214 35126 5323 35128
rect 5257 35123 5323 35126
rect 0 35050 800 35080
rect 1485 35050 1551 35053
rect 0 35048 1551 35050
rect 0 34992 1490 35048
rect 1546 34992 1551 35048
rect 0 34990 1551 34992
rect 0 34960 800 34990
rect 1485 34987 1551 34990
rect 4207 34848 4527 34849
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 34783 4527 34784
rect 7471 34848 7791 34849
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 34783 7791 34784
rect 10041 34642 10107 34645
rect 11200 34642 12000 34672
rect 10041 34640 12000 34642
rect 10041 34584 10046 34640
rect 10102 34584 12000 34640
rect 10041 34582 12000 34584
rect 10041 34579 10107 34582
rect 11200 34552 12000 34582
rect 0 34506 800 34536
rect 3049 34506 3115 34509
rect 0 34504 3115 34506
rect 0 34448 3054 34504
rect 3110 34448 3115 34504
rect 0 34446 3115 34448
rect 0 34416 800 34446
rect 3049 34443 3115 34446
rect 2576 34304 2896 34305
rect 2576 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2576 34239 2896 34240
rect 5839 34304 6159 34305
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 34239 6159 34240
rect 9103 34304 9423 34305
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 34239 9423 34240
rect 0 34098 800 34128
rect 3233 34098 3299 34101
rect 0 34096 3299 34098
rect 0 34040 3238 34096
rect 3294 34040 3299 34096
rect 0 34038 3299 34040
rect 0 34008 800 34038
rect 3233 34035 3299 34038
rect 2998 33764 3004 33828
rect 3068 33826 3074 33828
rect 3325 33826 3391 33829
rect 3068 33824 3391 33826
rect 3068 33768 3330 33824
rect 3386 33768 3391 33824
rect 3068 33766 3391 33768
rect 3068 33764 3074 33766
rect 3325 33763 3391 33766
rect 10041 33826 10107 33829
rect 11200 33826 12000 33856
rect 10041 33824 12000 33826
rect 10041 33768 10046 33824
rect 10102 33768 12000 33824
rect 10041 33766 12000 33768
rect 10041 33763 10107 33766
rect 4207 33760 4527 33761
rect 0 33690 800 33720
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 33695 4527 33696
rect 7471 33760 7791 33761
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 11200 33736 12000 33766
rect 7471 33695 7791 33696
rect 2313 33690 2379 33693
rect 0 33688 2379 33690
rect 0 33632 2318 33688
rect 2374 33632 2379 33688
rect 0 33630 2379 33632
rect 0 33600 800 33630
rect 2313 33627 2379 33630
rect 0 33282 800 33312
rect 1485 33282 1551 33285
rect 0 33280 1551 33282
rect 0 33224 1490 33280
rect 1546 33224 1551 33280
rect 0 33222 1551 33224
rect 0 33192 800 33222
rect 1485 33219 1551 33222
rect 2576 33216 2896 33217
rect 2576 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2576 33151 2896 33152
rect 5839 33216 6159 33217
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 33151 6159 33152
rect 9103 33216 9423 33217
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 33151 9423 33152
rect 10041 33010 10107 33013
rect 11200 33010 12000 33040
rect 10041 33008 12000 33010
rect 10041 32952 10046 33008
rect 10102 32952 12000 33008
rect 10041 32950 12000 32952
rect 10041 32947 10107 32950
rect 11200 32920 12000 32950
rect 0 32874 800 32904
rect 2313 32874 2379 32877
rect 0 32872 2379 32874
rect 0 32816 2318 32872
rect 2374 32816 2379 32872
rect 0 32814 2379 32816
rect 0 32784 800 32814
rect 2313 32811 2379 32814
rect 4207 32672 4527 32673
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 4207 32607 4527 32608
rect 7471 32672 7791 32673
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 32607 7791 32608
rect 2313 32604 2379 32605
rect 2262 32540 2268 32604
rect 2332 32602 2379 32604
rect 2332 32600 2424 32602
rect 2374 32544 2424 32600
rect 2332 32542 2424 32544
rect 2332 32540 2379 32542
rect 2313 32539 2379 32540
rect 0 32466 800 32496
rect 1393 32466 1459 32469
rect 0 32464 1459 32466
rect 0 32408 1398 32464
rect 1454 32408 1459 32464
rect 0 32406 1459 32408
rect 0 32376 800 32406
rect 1393 32403 1459 32406
rect 2078 32404 2084 32468
rect 2148 32466 2154 32468
rect 2497 32466 2563 32469
rect 2148 32464 2563 32466
rect 2148 32408 2502 32464
rect 2558 32408 2563 32464
rect 2148 32406 2563 32408
rect 2148 32404 2154 32406
rect 2497 32403 2563 32406
rect 10041 32330 10107 32333
rect 11200 32330 12000 32360
rect 10041 32328 12000 32330
rect 10041 32272 10046 32328
rect 10102 32272 12000 32328
rect 10041 32270 12000 32272
rect 10041 32267 10107 32270
rect 11200 32240 12000 32270
rect 2576 32128 2896 32129
rect 2576 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 2576 32063 2896 32064
rect 5839 32128 6159 32129
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 32063 6159 32064
rect 9103 32128 9423 32129
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 32063 9423 32064
rect 1526 31996 1532 32060
rect 1596 32058 1602 32060
rect 1669 32058 1735 32061
rect 1596 32056 1735 32058
rect 1596 32000 1674 32056
rect 1730 32000 1735 32056
rect 1596 31998 1735 32000
rect 1596 31996 1602 31998
rect 1669 31995 1735 31998
rect 0 31922 800 31952
rect 1209 31922 1275 31925
rect 0 31920 1275 31922
rect 0 31864 1214 31920
rect 1270 31864 1275 31920
rect 0 31862 1275 31864
rect 0 31832 800 31862
rect 1209 31859 1275 31862
rect 1761 31788 1827 31789
rect 1710 31724 1716 31788
rect 1780 31786 1827 31788
rect 1780 31784 1872 31786
rect 1822 31728 1872 31784
rect 1780 31726 1872 31728
rect 2221 31784 2287 31789
rect 2221 31728 2226 31784
rect 2282 31728 2287 31784
rect 1780 31724 1827 31726
rect 1761 31723 1827 31724
rect 2221 31723 2287 31728
rect 2224 31653 2284 31723
rect 2221 31648 2287 31653
rect 3601 31652 3667 31653
rect 3550 31650 3556 31652
rect 2221 31592 2226 31648
rect 2282 31592 2287 31648
rect 2221 31587 2287 31592
rect 3510 31590 3556 31650
rect 3620 31648 3667 31652
rect 3662 31592 3667 31648
rect 3550 31588 3556 31590
rect 3620 31588 3667 31592
rect 3601 31587 3667 31588
rect 4207 31584 4527 31585
rect 0 31514 800 31544
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 31519 4527 31520
rect 7471 31584 7791 31585
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 31519 7791 31520
rect 2405 31514 2471 31517
rect 0 31512 2471 31514
rect 0 31456 2410 31512
rect 2466 31456 2471 31512
rect 0 31454 2471 31456
rect 0 31424 800 31454
rect 2405 31451 2471 31454
rect 10041 31514 10107 31517
rect 11200 31514 12000 31544
rect 10041 31512 12000 31514
rect 10041 31456 10046 31512
rect 10102 31456 12000 31512
rect 10041 31454 12000 31456
rect 10041 31451 10107 31454
rect 11200 31424 12000 31454
rect 0 31106 800 31136
rect 2405 31106 2471 31109
rect 0 31104 2471 31106
rect 0 31048 2410 31104
rect 2466 31048 2471 31104
rect 0 31046 2471 31048
rect 0 31016 800 31046
rect 2405 31043 2471 31046
rect 2576 31040 2896 31041
rect 2576 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2576 30975 2896 30976
rect 5839 31040 6159 31041
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 30975 6159 30976
rect 9103 31040 9423 31041
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 30975 9423 30976
rect 10041 30834 10107 30837
rect 11200 30834 12000 30864
rect 10041 30832 12000 30834
rect 10041 30776 10046 30832
rect 10102 30776 12000 30832
rect 10041 30774 12000 30776
rect 10041 30771 10107 30774
rect 11200 30744 12000 30774
rect 0 30698 800 30728
rect 1485 30698 1551 30701
rect 0 30696 1551 30698
rect 0 30640 1490 30696
rect 1546 30640 1551 30696
rect 0 30638 1551 30640
rect 0 30608 800 30638
rect 1485 30635 1551 30638
rect 4207 30496 4527 30497
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 30431 4527 30432
rect 7471 30496 7791 30497
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 30431 7791 30432
rect 0 30290 800 30320
rect 2313 30290 2379 30293
rect 0 30288 2379 30290
rect 0 30232 2318 30288
rect 2374 30232 2379 30288
rect 0 30230 2379 30232
rect 0 30200 800 30230
rect 2313 30227 2379 30230
rect 10041 30018 10107 30021
rect 11200 30018 12000 30048
rect 10041 30016 12000 30018
rect 10041 29960 10046 30016
rect 10102 29960 12000 30016
rect 10041 29958 12000 29960
rect 10041 29955 10107 29958
rect 2576 29952 2896 29953
rect 0 29882 800 29912
rect 2576 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 2576 29887 2896 29888
rect 5839 29952 6159 29953
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 29887 6159 29888
rect 9103 29952 9423 29953
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 11200 29928 12000 29958
rect 9103 29887 9423 29888
rect 0 29822 1594 29882
rect 0 29792 800 29822
rect 1534 29746 1594 29822
rect 2957 29746 3023 29749
rect 1534 29744 3023 29746
rect 1534 29688 2962 29744
rect 3018 29688 3023 29744
rect 1534 29686 3023 29688
rect 2957 29683 3023 29686
rect 4207 29408 4527 29409
rect 0 29338 800 29368
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 4207 29343 4527 29344
rect 7471 29408 7791 29409
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 29343 7791 29344
rect 2129 29338 2195 29341
rect 0 29336 2195 29338
rect 0 29280 2134 29336
rect 2190 29280 2195 29336
rect 0 29278 2195 29280
rect 0 29248 800 29278
rect 2129 29275 2195 29278
rect 1761 29204 1827 29205
rect 1710 29202 1716 29204
rect 1670 29142 1716 29202
rect 1780 29200 1827 29204
rect 1822 29144 1827 29200
rect 1710 29140 1716 29142
rect 1780 29140 1827 29144
rect 1761 29139 1827 29140
rect 10961 29202 11027 29205
rect 11200 29202 12000 29232
rect 10961 29200 12000 29202
rect 10961 29144 10966 29200
rect 11022 29144 12000 29200
rect 10961 29142 12000 29144
rect 10961 29139 11027 29142
rect 11200 29112 12000 29142
rect 2773 29010 2839 29013
rect 2773 29008 3020 29010
rect 0 28930 800 28960
rect 2773 28952 2778 29008
rect 2834 28952 3020 29008
rect 2773 28950 3020 28952
rect 2773 28947 2839 28950
rect 2960 28932 3020 28950
rect 0 28870 1456 28930
rect 2960 28870 3004 28932
rect 0 28840 800 28870
rect 1396 28658 1456 28870
rect 2998 28868 3004 28870
rect 3068 28868 3074 28932
rect 2576 28864 2896 28865
rect 2576 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2576 28799 2896 28800
rect 5839 28864 6159 28865
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 28799 6159 28800
rect 9103 28864 9423 28865
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 28799 9423 28800
rect 3785 28658 3851 28661
rect 1396 28656 3851 28658
rect 1396 28600 3790 28656
rect 3846 28600 3851 28656
rect 1396 28598 3851 28600
rect 3785 28595 3851 28598
rect 0 28522 800 28552
rect 3417 28522 3483 28525
rect 0 28520 3483 28522
rect 0 28464 3422 28520
rect 3478 28464 3483 28520
rect 0 28462 3483 28464
rect 0 28432 800 28462
rect 3417 28459 3483 28462
rect 10133 28522 10199 28525
rect 11200 28522 12000 28552
rect 10133 28520 12000 28522
rect 10133 28464 10138 28520
rect 10194 28464 12000 28520
rect 10133 28462 12000 28464
rect 10133 28459 10199 28462
rect 11200 28432 12000 28462
rect 4207 28320 4527 28321
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 28255 4527 28256
rect 7471 28320 7791 28321
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 28255 7791 28256
rect 0 28114 800 28144
rect 1393 28114 1459 28117
rect 0 28112 1459 28114
rect 0 28056 1398 28112
rect 1454 28056 1459 28112
rect 0 28054 1459 28056
rect 0 28024 800 28054
rect 1393 28051 1459 28054
rect 3969 27978 4035 27981
rect 2086 27976 4035 27978
rect 2086 27920 3974 27976
rect 4030 27920 4035 27976
rect 2086 27918 4035 27920
rect 0 27706 800 27736
rect 2086 27706 2146 27918
rect 3969 27915 4035 27918
rect 2576 27776 2896 27777
rect 2576 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2576 27711 2896 27712
rect 5839 27776 6159 27777
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 27711 6159 27712
rect 9103 27776 9423 27777
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 27711 9423 27712
rect 0 27646 2146 27706
rect 10133 27706 10199 27709
rect 11200 27706 12000 27736
rect 10133 27704 12000 27706
rect 10133 27648 10138 27704
rect 10194 27648 12000 27704
rect 10133 27646 12000 27648
rect 0 27616 800 27646
rect 10133 27643 10199 27646
rect 11200 27616 12000 27646
rect 2773 27570 2839 27573
rect 3969 27570 4035 27573
rect 2773 27568 4035 27570
rect 2773 27512 2778 27568
rect 2834 27512 3974 27568
rect 4030 27512 4035 27568
rect 2773 27510 4035 27512
rect 2773 27507 2839 27510
rect 3969 27507 4035 27510
rect 2865 27434 2931 27437
rect 6269 27434 6335 27437
rect 2865 27432 6335 27434
rect 2865 27376 2870 27432
rect 2926 27376 6274 27432
rect 6330 27376 6335 27432
rect 2865 27374 6335 27376
rect 2865 27371 2931 27374
rect 6269 27371 6335 27374
rect 0 27298 800 27328
rect 3417 27298 3483 27301
rect 0 27296 3483 27298
rect 0 27240 3422 27296
rect 3478 27240 3483 27296
rect 0 27238 3483 27240
rect 0 27208 800 27238
rect 3417 27235 3483 27238
rect 4207 27232 4527 27233
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 4207 27167 4527 27168
rect 7471 27232 7791 27233
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 27167 7791 27168
rect 10133 27026 10199 27029
rect 11200 27026 12000 27056
rect 10133 27024 12000 27026
rect 10133 26968 10138 27024
rect 10194 26968 12000 27024
rect 10133 26966 12000 26968
rect 10133 26963 10199 26966
rect 11200 26936 12000 26966
rect 0 26890 800 26920
rect 3693 26890 3759 26893
rect 0 26888 3759 26890
rect 0 26832 3698 26888
rect 3754 26832 3759 26888
rect 0 26830 3759 26832
rect 0 26800 800 26830
rect 3693 26827 3759 26830
rect 2998 26692 3004 26756
rect 3068 26754 3074 26756
rect 3601 26754 3667 26757
rect 3068 26752 3667 26754
rect 3068 26696 3606 26752
rect 3662 26696 3667 26752
rect 3068 26694 3667 26696
rect 3068 26692 3074 26694
rect 3601 26691 3667 26694
rect 2576 26688 2896 26689
rect 2576 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2576 26623 2896 26624
rect 5839 26688 6159 26689
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 26623 6159 26624
rect 9103 26688 9423 26689
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 26623 9423 26624
rect 0 26346 800 26376
rect 3509 26346 3575 26349
rect 0 26344 3575 26346
rect 0 26288 3514 26344
rect 3570 26288 3575 26344
rect 0 26286 3575 26288
rect 0 26256 800 26286
rect 3509 26283 3575 26286
rect 10133 26210 10199 26213
rect 11200 26210 12000 26240
rect 10133 26208 12000 26210
rect 10133 26152 10138 26208
rect 10194 26152 12000 26208
rect 10133 26150 12000 26152
rect 10133 26147 10199 26150
rect 4207 26144 4527 26145
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 26079 4527 26080
rect 7471 26144 7791 26145
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 11200 26120 12000 26150
rect 7471 26079 7791 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 2129 25938 2195 25941
rect 2129 25936 2330 25938
rect 2129 25880 2134 25936
rect 2190 25880 2330 25936
rect 2129 25878 2330 25880
rect 2129 25875 2195 25878
rect 0 25530 800 25560
rect 1485 25530 1551 25533
rect 0 25528 1551 25530
rect 0 25472 1490 25528
rect 1546 25472 1551 25528
rect 0 25470 1551 25472
rect 0 25440 800 25470
rect 1485 25467 1551 25470
rect 2270 25394 2330 25878
rect 2576 25600 2896 25601
rect 2576 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2576 25535 2896 25536
rect 5839 25600 6159 25601
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 25535 6159 25536
rect 9103 25600 9423 25601
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 25535 9423 25536
rect 2589 25394 2655 25397
rect 2270 25392 2655 25394
rect 2270 25336 2594 25392
rect 2650 25336 2655 25392
rect 2270 25334 2655 25336
rect 2589 25331 2655 25334
rect 10225 25394 10291 25397
rect 11200 25394 12000 25424
rect 10225 25392 12000 25394
rect 10225 25336 10230 25392
rect 10286 25336 12000 25392
rect 10225 25334 12000 25336
rect 10225 25331 10291 25334
rect 11200 25304 12000 25334
rect 0 25122 800 25152
rect 2957 25122 3023 25125
rect 0 25120 3023 25122
rect 0 25064 2962 25120
rect 3018 25064 3023 25120
rect 0 25062 3023 25064
rect 0 25032 800 25062
rect 2957 25059 3023 25062
rect 4207 25056 4527 25057
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 24991 4527 24992
rect 7471 25056 7791 25057
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 24991 7791 24992
rect 0 24714 800 24744
rect 3233 24714 3299 24717
rect 0 24712 3299 24714
rect 0 24656 3238 24712
rect 3294 24656 3299 24712
rect 0 24654 3299 24656
rect 0 24624 800 24654
rect 3233 24651 3299 24654
rect 10133 24714 10199 24717
rect 11200 24714 12000 24744
rect 10133 24712 12000 24714
rect 10133 24656 10138 24712
rect 10194 24656 12000 24712
rect 10133 24654 12000 24656
rect 10133 24651 10199 24654
rect 11200 24624 12000 24654
rect 2576 24512 2896 24513
rect 2576 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2576 24447 2896 24448
rect 5839 24512 6159 24513
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 24447 6159 24448
rect 9103 24512 9423 24513
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 24447 9423 24448
rect 0 24306 800 24336
rect 1209 24306 1275 24309
rect 0 24304 1275 24306
rect 0 24248 1214 24304
rect 1270 24248 1275 24304
rect 0 24246 1275 24248
rect 0 24216 800 24246
rect 1209 24243 1275 24246
rect 4207 23968 4527 23969
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 23903 4527 23904
rect 7471 23968 7791 23969
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 23903 7791 23904
rect 10133 23898 10199 23901
rect 11200 23898 12000 23928
rect 10133 23896 12000 23898
rect 10133 23840 10138 23896
rect 10194 23840 12000 23896
rect 10133 23838 12000 23840
rect 10133 23835 10199 23838
rect 11200 23808 12000 23838
rect 0 23762 800 23792
rect 3141 23762 3207 23765
rect 0 23760 3207 23762
rect 0 23704 3146 23760
rect 3202 23704 3207 23760
rect 0 23702 3207 23704
rect 0 23672 800 23702
rect 3141 23699 3207 23702
rect 2576 23424 2896 23425
rect 0 23354 800 23384
rect 2576 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2576 23359 2896 23360
rect 5839 23424 6159 23425
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 23359 6159 23360
rect 9103 23424 9423 23425
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 23359 9423 23360
rect 1485 23354 1551 23357
rect 0 23352 1551 23354
rect 0 23296 1490 23352
rect 1546 23296 1551 23352
rect 0 23294 1551 23296
rect 0 23264 800 23294
rect 1485 23291 1551 23294
rect 10041 23218 10107 23221
rect 11200 23218 12000 23248
rect 10041 23216 12000 23218
rect 10041 23160 10046 23216
rect 10102 23160 12000 23216
rect 10041 23158 12000 23160
rect 10041 23155 10107 23158
rect 11200 23128 12000 23158
rect 0 22946 800 22976
rect 1393 22946 1459 22949
rect 0 22944 1459 22946
rect 0 22888 1398 22944
rect 1454 22888 1459 22944
rect 0 22886 1459 22888
rect 0 22856 800 22886
rect 1393 22883 1459 22886
rect 4207 22880 4527 22881
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 22815 4527 22816
rect 7471 22880 7791 22881
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 22815 7791 22816
rect 0 22538 800 22568
rect 3141 22538 3207 22541
rect 0 22536 3207 22538
rect 0 22480 3146 22536
rect 3202 22480 3207 22536
rect 0 22478 3207 22480
rect 0 22448 800 22478
rect 3141 22475 3207 22478
rect 10041 22402 10107 22405
rect 11200 22402 12000 22432
rect 10041 22400 12000 22402
rect 10041 22344 10046 22400
rect 10102 22344 12000 22400
rect 10041 22342 12000 22344
rect 10041 22339 10107 22342
rect 2576 22336 2896 22337
rect 2576 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2576 22271 2896 22272
rect 5839 22336 6159 22337
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 22271 6159 22272
rect 9103 22336 9423 22337
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 11200 22312 12000 22342
rect 9103 22271 9423 22272
rect 0 22130 800 22160
rect 1209 22130 1275 22133
rect 0 22128 1275 22130
rect 0 22072 1214 22128
rect 1270 22072 1275 22128
rect 0 22070 1275 22072
rect 0 22040 800 22070
rect 1209 22067 1275 22070
rect 4207 21792 4527 21793
rect 0 21722 800 21752
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 21727 4527 21728
rect 7471 21792 7791 21793
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 21727 7791 21728
rect 3969 21722 4035 21725
rect 0 21720 4035 21722
rect 0 21664 3974 21720
rect 4030 21664 4035 21720
rect 0 21662 4035 21664
rect 0 21632 800 21662
rect 3969 21659 4035 21662
rect 10041 21586 10107 21589
rect 11200 21586 12000 21616
rect 10041 21584 12000 21586
rect 10041 21528 10046 21584
rect 10102 21528 12000 21584
rect 10041 21526 12000 21528
rect 10041 21523 10107 21526
rect 11200 21496 12000 21526
rect 2865 21450 2931 21453
rect 1396 21448 2931 21450
rect 1396 21392 2870 21448
rect 2926 21392 2931 21448
rect 1396 21390 2931 21392
rect 0 21178 800 21208
rect 1396 21178 1456 21390
rect 2865 21387 2931 21390
rect 2576 21248 2896 21249
rect 2576 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2576 21183 2896 21184
rect 5839 21248 6159 21249
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 21183 6159 21184
rect 9103 21248 9423 21249
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 21183 9423 21184
rect 0 21118 1456 21178
rect 0 21088 800 21118
rect 10041 20906 10107 20909
rect 11200 20906 12000 20936
rect 10041 20904 12000 20906
rect 10041 20848 10046 20904
rect 10102 20848 12000 20904
rect 10041 20846 12000 20848
rect 10041 20843 10107 20846
rect 11200 20816 12000 20846
rect 0 20770 800 20800
rect 3877 20770 3943 20773
rect 0 20768 3943 20770
rect 0 20712 3882 20768
rect 3938 20712 3943 20768
rect 0 20710 3943 20712
rect 0 20680 800 20710
rect 3877 20707 3943 20710
rect 4207 20704 4527 20705
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 20639 4527 20640
rect 7471 20704 7791 20705
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 20639 7791 20640
rect 0 20362 800 20392
rect 3969 20362 4035 20365
rect 0 20360 4035 20362
rect 0 20304 3974 20360
rect 4030 20304 4035 20360
rect 0 20302 4035 20304
rect 0 20272 800 20302
rect 3969 20299 4035 20302
rect 2576 20160 2896 20161
rect 2576 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2576 20095 2896 20096
rect 5839 20160 6159 20161
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 20095 6159 20096
rect 9103 20160 9423 20161
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 20095 9423 20096
rect 10041 20090 10107 20093
rect 11200 20090 12000 20120
rect 10041 20088 12000 20090
rect 10041 20032 10046 20088
rect 10102 20032 12000 20088
rect 10041 20030 12000 20032
rect 10041 20027 10107 20030
rect 11200 20000 12000 20030
rect 0 19954 800 19984
rect 4061 19954 4127 19957
rect 0 19952 4127 19954
rect 0 19896 4066 19952
rect 4122 19896 4127 19952
rect 0 19894 4127 19896
rect 0 19864 800 19894
rect 4061 19891 4127 19894
rect 4207 19616 4527 19617
rect 0 19546 800 19576
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 19551 4527 19552
rect 7471 19616 7791 19617
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 19551 7791 19552
rect 3417 19546 3483 19549
rect 0 19544 3483 19546
rect 0 19488 3422 19544
rect 3478 19488 3483 19544
rect 0 19486 3483 19488
rect 0 19456 800 19486
rect 3417 19483 3483 19486
rect 10041 19410 10107 19413
rect 11200 19410 12000 19440
rect 10041 19408 12000 19410
rect 10041 19352 10046 19408
rect 10102 19352 12000 19408
rect 10041 19350 12000 19352
rect 10041 19347 10107 19350
rect 11200 19320 12000 19350
rect 3049 19274 3115 19277
rect 1396 19272 3115 19274
rect 1396 19216 3054 19272
rect 3110 19216 3115 19272
rect 1396 19214 3115 19216
rect 0 19138 800 19168
rect 1396 19138 1456 19214
rect 3049 19211 3115 19214
rect 0 19078 1456 19138
rect 0 19048 800 19078
rect 2576 19072 2896 19073
rect 2576 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2576 19007 2896 19008
rect 5839 19072 6159 19073
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 19007 6159 19008
rect 9103 19072 9423 19073
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 19007 9423 19008
rect 0 18594 800 18624
rect 3233 18594 3299 18597
rect 0 18592 3299 18594
rect 0 18536 3238 18592
rect 3294 18536 3299 18592
rect 0 18534 3299 18536
rect 0 18504 800 18534
rect 3233 18531 3299 18534
rect 10041 18594 10107 18597
rect 11200 18594 12000 18624
rect 10041 18592 12000 18594
rect 10041 18536 10046 18592
rect 10102 18536 12000 18592
rect 10041 18534 12000 18536
rect 10041 18531 10107 18534
rect 4207 18528 4527 18529
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 18463 4527 18464
rect 7471 18528 7791 18529
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 11200 18504 12000 18534
rect 7471 18463 7791 18464
rect 0 18186 800 18216
rect 2773 18186 2839 18189
rect 0 18184 2839 18186
rect 0 18128 2778 18184
rect 2834 18128 2839 18184
rect 0 18126 2839 18128
rect 0 18096 800 18126
rect 2773 18123 2839 18126
rect 2576 17984 2896 17985
rect 2576 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2576 17919 2896 17920
rect 5839 17984 6159 17985
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 17919 6159 17920
rect 9103 17984 9423 17985
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 17919 9423 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 10041 17778 10107 17781
rect 11200 17778 12000 17808
rect 10041 17776 12000 17778
rect 10041 17720 10046 17776
rect 10102 17720 12000 17776
rect 10041 17718 12000 17720
rect 10041 17715 10107 17718
rect 11200 17688 12000 17718
rect 4207 17440 4527 17441
rect 0 17370 800 17400
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 17375 4527 17376
rect 7471 17440 7791 17441
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 17375 7791 17376
rect 3049 17370 3115 17373
rect 0 17368 3115 17370
rect 0 17312 3054 17368
rect 3110 17312 3115 17368
rect 0 17310 3115 17312
rect 0 17280 800 17310
rect 3049 17307 3115 17310
rect 2865 17098 2931 17101
rect 1396 17096 2931 17098
rect 1396 17040 2870 17096
rect 2926 17040 2931 17096
rect 1396 17038 2931 17040
rect 0 16962 800 16992
rect 1396 16962 1456 17038
rect 2865 17035 2931 17038
rect 10041 17098 10107 17101
rect 11200 17098 12000 17128
rect 10041 17096 12000 17098
rect 10041 17040 10046 17096
rect 10102 17040 12000 17096
rect 10041 17038 12000 17040
rect 10041 17035 10107 17038
rect 11200 17008 12000 17038
rect 0 16902 1456 16962
rect 0 16872 800 16902
rect 2576 16896 2896 16897
rect 2576 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2576 16831 2896 16832
rect 5839 16896 6159 16897
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 16831 6159 16832
rect 9103 16896 9423 16897
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 16831 9423 16832
rect 0 16554 800 16584
rect 2221 16554 2287 16557
rect 0 16552 2287 16554
rect 0 16496 2226 16552
rect 2282 16496 2287 16552
rect 0 16494 2287 16496
rect 0 16464 800 16494
rect 2221 16491 2287 16494
rect 4207 16352 4527 16353
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 16287 4527 16288
rect 7471 16352 7791 16353
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 16287 7791 16288
rect 10041 16282 10107 16285
rect 11200 16282 12000 16312
rect 10041 16280 12000 16282
rect 10041 16224 10046 16280
rect 10102 16224 12000 16280
rect 10041 16222 12000 16224
rect 10041 16219 10107 16222
rect 11200 16192 12000 16222
rect 0 16010 800 16040
rect 3233 16010 3299 16013
rect 0 16008 3299 16010
rect 0 15952 3238 16008
rect 3294 15952 3299 16008
rect 0 15950 3299 15952
rect 0 15920 800 15950
rect 3233 15947 3299 15950
rect 2576 15808 2896 15809
rect 2576 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2576 15743 2896 15744
rect 5839 15808 6159 15809
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 15743 6159 15744
rect 9103 15808 9423 15809
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 15743 9423 15744
rect 0 15602 800 15632
rect 1209 15602 1275 15605
rect 0 15600 1275 15602
rect 0 15544 1214 15600
rect 1270 15544 1275 15600
rect 0 15542 1275 15544
rect 0 15512 800 15542
rect 1209 15539 1275 15542
rect 10041 15602 10107 15605
rect 11200 15602 12000 15632
rect 10041 15600 12000 15602
rect 10041 15544 10046 15600
rect 10102 15544 12000 15600
rect 10041 15542 12000 15544
rect 10041 15539 10107 15542
rect 11200 15512 12000 15542
rect 4207 15264 4527 15265
rect 0 15194 800 15224
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 15199 4527 15200
rect 7471 15264 7791 15265
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 15199 7791 15200
rect 1853 15194 1919 15197
rect 0 15192 1919 15194
rect 0 15136 1858 15192
rect 1914 15136 1919 15192
rect 0 15134 1919 15136
rect 0 15104 800 15134
rect 1853 15131 1919 15134
rect 2773 15194 2839 15197
rect 3601 15194 3667 15197
rect 2773 15192 3667 15194
rect 2773 15136 2778 15192
rect 2834 15136 3606 15192
rect 3662 15136 3667 15192
rect 2773 15134 3667 15136
rect 2773 15131 2839 15134
rect 3601 15131 3667 15134
rect 3233 14922 3299 14925
rect 3877 14922 3943 14925
rect 3233 14920 3943 14922
rect 3233 14864 3238 14920
rect 3294 14864 3882 14920
rect 3938 14864 3943 14920
rect 3233 14862 3943 14864
rect 3233 14859 3299 14862
rect 3877 14859 3943 14862
rect 0 14786 800 14816
rect 1117 14786 1183 14789
rect 0 14784 1183 14786
rect 0 14728 1122 14784
rect 1178 14728 1183 14784
rect 0 14726 1183 14728
rect 0 14696 800 14726
rect 1117 14723 1183 14726
rect 10041 14786 10107 14789
rect 11200 14786 12000 14816
rect 10041 14784 12000 14786
rect 10041 14728 10046 14784
rect 10102 14728 12000 14784
rect 10041 14726 12000 14728
rect 10041 14723 10107 14726
rect 2576 14720 2896 14721
rect 2576 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2576 14655 2896 14656
rect 5839 14720 6159 14721
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 14655 6159 14656
rect 9103 14720 9423 14721
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 11200 14696 12000 14726
rect 9103 14655 9423 14656
rect 0 14378 800 14408
rect 4153 14378 4219 14381
rect 0 14376 4219 14378
rect 0 14320 4158 14376
rect 4214 14320 4219 14376
rect 0 14318 4219 14320
rect 0 14288 800 14318
rect 4153 14315 4219 14318
rect 4207 14176 4527 14177
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 14111 4527 14112
rect 7471 14176 7791 14177
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 14111 7791 14112
rect 0 13970 800 14000
rect 3969 13970 4035 13973
rect 0 13968 4035 13970
rect 0 13912 3974 13968
rect 4030 13912 4035 13968
rect 0 13910 4035 13912
rect 0 13880 800 13910
rect 3969 13907 4035 13910
rect 10041 13970 10107 13973
rect 11200 13970 12000 14000
rect 10041 13968 12000 13970
rect 10041 13912 10046 13968
rect 10102 13912 12000 13968
rect 10041 13910 12000 13912
rect 10041 13907 10107 13910
rect 11200 13880 12000 13910
rect 2576 13632 2896 13633
rect 0 13562 800 13592
rect 2576 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2576 13567 2896 13568
rect 5839 13632 6159 13633
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 13567 6159 13568
rect 9103 13632 9423 13633
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 13567 9423 13568
rect 0 13502 1456 13562
rect 0 13472 800 13502
rect 1396 13426 1456 13502
rect 4061 13426 4127 13429
rect 1396 13424 4127 13426
rect 1396 13368 4066 13424
rect 4122 13368 4127 13424
rect 1396 13366 4127 13368
rect 4061 13363 4127 13366
rect 10041 13290 10107 13293
rect 11200 13290 12000 13320
rect 10041 13288 12000 13290
rect 10041 13232 10046 13288
rect 10102 13232 12000 13288
rect 10041 13230 12000 13232
rect 10041 13227 10107 13230
rect 11200 13200 12000 13230
rect 4207 13088 4527 13089
rect 0 13018 800 13048
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 13023 4527 13024
rect 7471 13088 7791 13089
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 13023 7791 13024
rect 1853 13018 1919 13021
rect 0 13016 1919 13018
rect 0 12960 1858 13016
rect 1914 12960 1919 13016
rect 0 12958 1919 12960
rect 0 12928 800 12958
rect 1853 12955 1919 12958
rect 2773 12746 2839 12749
rect 1396 12744 2839 12746
rect 1396 12688 2778 12744
rect 2834 12688 2839 12744
rect 1396 12686 2839 12688
rect 0 12610 800 12640
rect 1396 12610 1456 12686
rect 2773 12683 2839 12686
rect 0 12550 1456 12610
rect 0 12520 800 12550
rect 2576 12544 2896 12545
rect 2576 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2576 12479 2896 12480
rect 5839 12544 6159 12545
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 12479 6159 12480
rect 9103 12544 9423 12545
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 12479 9423 12480
rect 10041 12474 10107 12477
rect 11200 12474 12000 12504
rect 10041 12472 12000 12474
rect 10041 12416 10046 12472
rect 10102 12416 12000 12472
rect 10041 12414 12000 12416
rect 10041 12411 10107 12414
rect 11200 12384 12000 12414
rect 1393 12338 1459 12341
rect 798 12336 1459 12338
rect 798 12280 1398 12336
rect 1454 12280 1459 12336
rect 798 12278 1459 12280
rect 798 12232 858 12278
rect 1393 12275 1459 12278
rect 0 12142 858 12232
rect 0 12112 800 12142
rect 4207 12000 4527 12001
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 11935 4527 11936
rect 7471 12000 7791 12001
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 11935 7791 11936
rect 0 11794 800 11824
rect 1485 11794 1551 11797
rect 0 11792 1551 11794
rect 0 11736 1490 11792
rect 1546 11736 1551 11792
rect 0 11734 1551 11736
rect 0 11704 800 11734
rect 1485 11731 1551 11734
rect 10041 11794 10107 11797
rect 11200 11794 12000 11824
rect 10041 11792 12000 11794
rect 10041 11736 10046 11792
rect 10102 11736 12000 11792
rect 10041 11734 12000 11736
rect 10041 11731 10107 11734
rect 11200 11704 12000 11734
rect 2576 11456 2896 11457
rect 0 11386 800 11416
rect 2576 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2576 11391 2896 11392
rect 5839 11456 6159 11457
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 11391 6159 11392
rect 9103 11456 9423 11457
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 11391 9423 11392
rect 1393 11386 1459 11389
rect 0 11384 1459 11386
rect 0 11328 1398 11384
rect 1454 11328 1459 11384
rect 0 11326 1459 11328
rect 0 11296 800 11326
rect 1393 11323 1459 11326
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 10041 10978 10107 10981
rect 11200 10978 12000 11008
rect 10041 10976 12000 10978
rect 10041 10920 10046 10976
rect 10102 10920 12000 10976
rect 10041 10918 12000 10920
rect 10041 10915 10107 10918
rect 4207 10912 4527 10913
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 10847 4527 10848
rect 7471 10912 7791 10913
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 11200 10888 12000 10918
rect 7471 10847 7791 10848
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 2576 10368 2896 10369
rect 2576 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2576 10303 2896 10304
rect 5839 10368 6159 10369
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 10303 6159 10304
rect 9103 10368 9423 10369
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 10303 9423 10304
rect 10041 10162 10107 10165
rect 11200 10162 12000 10192
rect 10041 10160 12000 10162
rect 10041 10104 10046 10160
rect 10102 10104 12000 10160
rect 10041 10102 12000 10104
rect 10041 10099 10107 10102
rect 11200 10072 12000 10102
rect 0 10026 800 10056
rect 1301 10026 1367 10029
rect 0 10024 1367 10026
rect 0 9968 1306 10024
rect 1362 9968 1367 10024
rect 0 9966 1367 9968
rect 0 9936 800 9966
rect 1301 9963 1367 9966
rect 4207 9824 4527 9825
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 9759 4527 9760
rect 7471 9824 7791 9825
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 9759 7791 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 10041 9482 10107 9485
rect 11200 9482 12000 9512
rect 10041 9480 12000 9482
rect 10041 9424 10046 9480
rect 10102 9424 12000 9480
rect 10041 9422 12000 9424
rect 10041 9419 10107 9422
rect 11200 9392 12000 9422
rect 2576 9280 2896 9281
rect 0 9210 800 9240
rect 2576 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2576 9215 2896 9216
rect 5839 9280 6159 9281
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 9215 6159 9216
rect 9103 9280 9423 9281
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 9215 9423 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 0 8802 800 8832
rect 3785 8802 3851 8805
rect 0 8800 3851 8802
rect 0 8744 3790 8800
rect 3846 8744 3851 8800
rect 0 8742 3851 8744
rect 0 8712 800 8742
rect 3785 8739 3851 8742
rect 4207 8736 4527 8737
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 8671 4527 8672
rect 7471 8736 7791 8737
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 8671 7791 8672
rect 10041 8666 10107 8669
rect 11200 8666 12000 8696
rect 10041 8664 12000 8666
rect 10041 8608 10046 8664
rect 10102 8608 12000 8664
rect 10041 8606 12000 8608
rect 10041 8603 10107 8606
rect 11200 8576 12000 8606
rect 0 8394 800 8424
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 2576 8192 2896 8193
rect 2576 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2576 8127 2896 8128
rect 5839 8192 6159 8193
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 8127 6159 8128
rect 9103 8192 9423 8193
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 8127 9423 8128
rect 10041 7986 10107 7989
rect 11200 7986 12000 8016
rect 10041 7984 12000 7986
rect 10041 7928 10046 7984
rect 10102 7928 12000 7984
rect 10041 7926 12000 7928
rect 10041 7923 10107 7926
rect 11200 7896 12000 7926
rect 0 7850 800 7880
rect 1301 7850 1367 7853
rect 0 7848 1367 7850
rect 0 7792 1306 7848
rect 1362 7792 1367 7848
rect 0 7790 1367 7792
rect 0 7760 800 7790
rect 1301 7787 1367 7790
rect 4207 7648 4527 7649
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 7583 4527 7584
rect 7471 7648 7791 7649
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 7583 7791 7584
rect 0 7442 800 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 800 7382
rect 1393 7379 1459 7382
rect 2773 7306 2839 7309
rect 1350 7304 2839 7306
rect 1350 7248 2778 7304
rect 2834 7248 2839 7304
rect 1350 7246 2839 7248
rect 0 7034 800 7064
rect 1350 7034 1410 7246
rect 2773 7243 2839 7246
rect 10041 7170 10107 7173
rect 11200 7170 12000 7200
rect 10041 7168 12000 7170
rect 10041 7112 10046 7168
rect 10102 7112 12000 7168
rect 10041 7110 12000 7112
rect 10041 7107 10107 7110
rect 2576 7104 2896 7105
rect 2576 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2576 7039 2896 7040
rect 5839 7104 6159 7105
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 7039 6159 7040
rect 9103 7104 9423 7105
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 11200 7080 12000 7110
rect 9103 7039 9423 7040
rect 0 6974 1410 7034
rect 0 6944 800 6974
rect 0 6626 800 6656
rect 1853 6626 1919 6629
rect 0 6624 1919 6626
rect 0 6568 1858 6624
rect 1914 6568 1919 6624
rect 0 6566 1919 6568
rect 0 6536 800 6566
rect 1853 6563 1919 6566
rect 4207 6560 4527 6561
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 6495 4527 6496
rect 7471 6560 7791 6561
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 6495 7791 6496
rect 10041 6354 10107 6357
rect 11200 6354 12000 6384
rect 10041 6352 12000 6354
rect 10041 6296 10046 6352
rect 10102 6296 12000 6352
rect 10041 6294 12000 6296
rect 10041 6291 10107 6294
rect 11200 6264 12000 6294
rect 0 6218 800 6248
rect 3785 6218 3851 6221
rect 0 6216 3851 6218
rect 0 6160 3790 6216
rect 3846 6160 3851 6216
rect 0 6158 3851 6160
rect 0 6128 800 6158
rect 3785 6155 3851 6158
rect 2576 6016 2896 6017
rect 2576 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2576 5951 2896 5952
rect 5839 6016 6159 6017
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 5951 6159 5952
rect 9103 6016 9423 6017
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 5951 9423 5952
rect 0 5810 800 5840
rect 3417 5810 3483 5813
rect 0 5808 3483 5810
rect 0 5752 3422 5808
rect 3478 5752 3483 5808
rect 0 5750 3483 5752
rect 0 5720 800 5750
rect 3417 5747 3483 5750
rect 10041 5674 10107 5677
rect 11200 5674 12000 5704
rect 10041 5672 12000 5674
rect 10041 5616 10046 5672
rect 10102 5616 12000 5672
rect 10041 5614 12000 5616
rect 10041 5611 10107 5614
rect 11200 5584 12000 5614
rect 4207 5472 4527 5473
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 5407 4527 5408
rect 7471 5472 7791 5473
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 5407 7791 5408
rect 0 5266 800 5296
rect 3969 5266 4035 5269
rect 0 5264 4035 5266
rect 0 5208 3974 5264
rect 4030 5208 4035 5264
rect 0 5206 4035 5208
rect 0 5176 800 5206
rect 3969 5203 4035 5206
rect 2576 4928 2896 4929
rect 0 4858 800 4888
rect 2576 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2576 4863 2896 4864
rect 5839 4928 6159 4929
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 4863 6159 4864
rect 9103 4928 9423 4929
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 4863 9423 4864
rect 10041 4858 10107 4861
rect 11200 4858 12000 4888
rect 0 4798 1594 4858
rect 0 4768 800 4798
rect 1534 4722 1594 4798
rect 10041 4856 12000 4858
rect 10041 4800 10046 4856
rect 10102 4800 12000 4856
rect 10041 4798 12000 4800
rect 10041 4795 10107 4798
rect 11200 4768 12000 4798
rect 2957 4722 3023 4725
rect 1534 4720 3023 4722
rect 1534 4664 2962 4720
rect 3018 4664 3023 4720
rect 1534 4662 3023 4664
rect 2957 4659 3023 4662
rect 0 4450 800 4480
rect 3969 4450 4035 4453
rect 0 4448 4035 4450
rect 0 4392 3974 4448
rect 4030 4392 4035 4448
rect 0 4390 4035 4392
rect 0 4360 800 4390
rect 3969 4387 4035 4390
rect 4207 4384 4527 4385
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 4319 4527 4320
rect 7471 4384 7791 4385
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 4319 7791 4320
rect 10041 4178 10107 4181
rect 11200 4178 12000 4208
rect 10041 4176 12000 4178
rect 10041 4120 10046 4176
rect 10102 4120 12000 4176
rect 10041 4118 12000 4120
rect 10041 4115 10107 4118
rect 11200 4088 12000 4118
rect 0 4042 800 4072
rect 3601 4042 3667 4045
rect 0 4040 3667 4042
rect 0 3984 3606 4040
rect 3662 3984 3667 4040
rect 0 3982 3667 3984
rect 0 3952 800 3982
rect 3601 3979 3667 3982
rect 2576 3840 2896 3841
rect 2576 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2576 3775 2896 3776
rect 5839 3840 6159 3841
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 3775 6159 3776
rect 9103 3840 9423 3841
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 3775 9423 3776
rect 0 3634 800 3664
rect 2865 3634 2931 3637
rect 0 3632 2931 3634
rect 0 3576 2870 3632
rect 2926 3576 2931 3632
rect 0 3574 2931 3576
rect 0 3544 800 3574
rect 2865 3571 2931 3574
rect 10041 3362 10107 3365
rect 11200 3362 12000 3392
rect 10041 3360 12000 3362
rect 10041 3304 10046 3360
rect 10102 3304 12000 3360
rect 10041 3302 12000 3304
rect 10041 3299 10107 3302
rect 4207 3296 4527 3297
rect 0 3226 800 3256
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 3231 4527 3232
rect 7471 3296 7791 3297
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 11200 3272 12000 3302
rect 7471 3231 7791 3232
rect 1301 3226 1367 3229
rect 0 3224 1367 3226
rect 0 3168 1306 3224
rect 1362 3168 1367 3224
rect 0 3166 1367 3168
rect 0 3136 800 3166
rect 1301 3163 1367 3166
rect 2576 2752 2896 2753
rect 0 2682 800 2712
rect 2576 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2576 2687 2896 2688
rect 5839 2752 6159 2753
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2687 6159 2688
rect 9103 2752 9423 2753
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2687 9423 2688
rect 1393 2682 1459 2685
rect 0 2680 1459 2682
rect 0 2624 1398 2680
rect 1454 2624 1459 2680
rect 0 2622 1459 2624
rect 0 2592 800 2622
rect 1393 2619 1459 2622
rect 10041 2546 10107 2549
rect 11200 2546 12000 2576
rect 10041 2544 12000 2546
rect 10041 2488 10046 2544
rect 10102 2488 12000 2544
rect 10041 2486 12000 2488
rect 10041 2483 10107 2486
rect 11200 2456 12000 2486
rect 0 2274 800 2304
rect 3509 2274 3575 2277
rect 0 2272 3575 2274
rect 0 2216 3514 2272
rect 3570 2216 3575 2272
rect 0 2214 3575 2216
rect 0 2184 800 2214
rect 3509 2211 3575 2214
rect 4207 2208 4527 2209
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2143 4527 2144
rect 7471 2208 7791 2209
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2143 7791 2144
rect 0 1866 800 1896
rect 3969 1866 4035 1869
rect 0 1864 4035 1866
rect 0 1808 3974 1864
rect 4030 1808 4035 1864
rect 0 1806 4035 1808
rect 0 1776 800 1806
rect 3969 1803 4035 1806
rect 9489 1866 9555 1869
rect 11200 1866 12000 1896
rect 9489 1864 12000 1866
rect 9489 1808 9494 1864
rect 9550 1808 12000 1864
rect 9489 1806 12000 1808
rect 9489 1803 9555 1806
rect 11200 1776 12000 1806
rect 0 1458 800 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 800 1398
rect 2865 1395 2931 1398
rect 0 1050 800 1080
rect 3601 1050 3667 1053
rect 0 1048 3667 1050
rect 0 992 3606 1048
rect 3662 992 3667 1048
rect 0 990 3667 992
rect 0 960 800 990
rect 3601 987 3667 990
rect 10041 1050 10107 1053
rect 11200 1050 12000 1080
rect 10041 1048 12000 1050
rect 10041 992 10046 1048
rect 10102 992 12000 1048
rect 10041 990 12000 992
rect 10041 987 10107 990
rect 11200 960 12000 990
rect 0 642 800 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 800 582
rect 2773 579 2839 582
rect 9305 370 9371 373
rect 11200 370 12000 400
rect 9305 368 12000 370
rect 9305 312 9310 368
rect 9366 312 12000 368
rect 9305 310 12000 312
rect 9305 307 9371 310
rect 11200 280 12000 310
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
<< via3 >>
rect 2584 77820 2648 77824
rect 2584 77764 2588 77820
rect 2588 77764 2644 77820
rect 2644 77764 2648 77820
rect 2584 77760 2648 77764
rect 2664 77820 2728 77824
rect 2664 77764 2668 77820
rect 2668 77764 2724 77820
rect 2724 77764 2728 77820
rect 2664 77760 2728 77764
rect 2744 77820 2808 77824
rect 2744 77764 2748 77820
rect 2748 77764 2804 77820
rect 2804 77764 2808 77820
rect 2744 77760 2808 77764
rect 2824 77820 2888 77824
rect 2824 77764 2828 77820
rect 2828 77764 2884 77820
rect 2884 77764 2888 77820
rect 2824 77760 2888 77764
rect 5847 77820 5911 77824
rect 5847 77764 5851 77820
rect 5851 77764 5907 77820
rect 5907 77764 5911 77820
rect 5847 77760 5911 77764
rect 5927 77820 5991 77824
rect 5927 77764 5931 77820
rect 5931 77764 5987 77820
rect 5987 77764 5991 77820
rect 5927 77760 5991 77764
rect 6007 77820 6071 77824
rect 6007 77764 6011 77820
rect 6011 77764 6067 77820
rect 6067 77764 6071 77820
rect 6007 77760 6071 77764
rect 6087 77820 6151 77824
rect 6087 77764 6091 77820
rect 6091 77764 6147 77820
rect 6147 77764 6151 77820
rect 6087 77760 6151 77764
rect 9111 77820 9175 77824
rect 9111 77764 9115 77820
rect 9115 77764 9171 77820
rect 9171 77764 9175 77820
rect 9111 77760 9175 77764
rect 9191 77820 9255 77824
rect 9191 77764 9195 77820
rect 9195 77764 9251 77820
rect 9251 77764 9255 77820
rect 9191 77760 9255 77764
rect 9271 77820 9335 77824
rect 9271 77764 9275 77820
rect 9275 77764 9331 77820
rect 9331 77764 9335 77820
rect 9271 77760 9335 77764
rect 9351 77820 9415 77824
rect 9351 77764 9355 77820
rect 9355 77764 9411 77820
rect 9411 77764 9415 77820
rect 9351 77760 9415 77764
rect 4215 77276 4279 77280
rect 4215 77220 4219 77276
rect 4219 77220 4275 77276
rect 4275 77220 4279 77276
rect 4215 77216 4279 77220
rect 4295 77276 4359 77280
rect 4295 77220 4299 77276
rect 4299 77220 4355 77276
rect 4355 77220 4359 77276
rect 4295 77216 4359 77220
rect 4375 77276 4439 77280
rect 4375 77220 4379 77276
rect 4379 77220 4435 77276
rect 4435 77220 4439 77276
rect 4375 77216 4439 77220
rect 4455 77276 4519 77280
rect 4455 77220 4459 77276
rect 4459 77220 4515 77276
rect 4515 77220 4519 77276
rect 4455 77216 4519 77220
rect 7479 77276 7543 77280
rect 7479 77220 7483 77276
rect 7483 77220 7539 77276
rect 7539 77220 7543 77276
rect 7479 77216 7543 77220
rect 7559 77276 7623 77280
rect 7559 77220 7563 77276
rect 7563 77220 7619 77276
rect 7619 77220 7623 77276
rect 7559 77216 7623 77220
rect 7639 77276 7703 77280
rect 7639 77220 7643 77276
rect 7643 77220 7699 77276
rect 7699 77220 7703 77276
rect 7639 77216 7703 77220
rect 7719 77276 7783 77280
rect 7719 77220 7723 77276
rect 7723 77220 7779 77276
rect 7779 77220 7783 77276
rect 7719 77216 7783 77220
rect 2584 76732 2648 76736
rect 2584 76676 2588 76732
rect 2588 76676 2644 76732
rect 2644 76676 2648 76732
rect 2584 76672 2648 76676
rect 2664 76732 2728 76736
rect 2664 76676 2668 76732
rect 2668 76676 2724 76732
rect 2724 76676 2728 76732
rect 2664 76672 2728 76676
rect 2744 76732 2808 76736
rect 2744 76676 2748 76732
rect 2748 76676 2804 76732
rect 2804 76676 2808 76732
rect 2744 76672 2808 76676
rect 2824 76732 2888 76736
rect 2824 76676 2828 76732
rect 2828 76676 2884 76732
rect 2884 76676 2888 76732
rect 2824 76672 2888 76676
rect 5847 76732 5911 76736
rect 5847 76676 5851 76732
rect 5851 76676 5907 76732
rect 5907 76676 5911 76732
rect 5847 76672 5911 76676
rect 5927 76732 5991 76736
rect 5927 76676 5931 76732
rect 5931 76676 5987 76732
rect 5987 76676 5991 76732
rect 5927 76672 5991 76676
rect 6007 76732 6071 76736
rect 6007 76676 6011 76732
rect 6011 76676 6067 76732
rect 6067 76676 6071 76732
rect 6007 76672 6071 76676
rect 6087 76732 6151 76736
rect 6087 76676 6091 76732
rect 6091 76676 6147 76732
rect 6147 76676 6151 76732
rect 6087 76672 6151 76676
rect 9111 76732 9175 76736
rect 9111 76676 9115 76732
rect 9115 76676 9171 76732
rect 9171 76676 9175 76732
rect 9111 76672 9175 76676
rect 9191 76732 9255 76736
rect 9191 76676 9195 76732
rect 9195 76676 9251 76732
rect 9251 76676 9255 76732
rect 9191 76672 9255 76676
rect 9271 76732 9335 76736
rect 9271 76676 9275 76732
rect 9275 76676 9331 76732
rect 9331 76676 9335 76732
rect 9271 76672 9335 76676
rect 9351 76732 9415 76736
rect 9351 76676 9355 76732
rect 9355 76676 9411 76732
rect 9411 76676 9415 76732
rect 9351 76672 9415 76676
rect 4215 76188 4279 76192
rect 4215 76132 4219 76188
rect 4219 76132 4275 76188
rect 4275 76132 4279 76188
rect 4215 76128 4279 76132
rect 4295 76188 4359 76192
rect 4295 76132 4299 76188
rect 4299 76132 4355 76188
rect 4355 76132 4359 76188
rect 4295 76128 4359 76132
rect 4375 76188 4439 76192
rect 4375 76132 4379 76188
rect 4379 76132 4435 76188
rect 4435 76132 4439 76188
rect 4375 76128 4439 76132
rect 4455 76188 4519 76192
rect 4455 76132 4459 76188
rect 4459 76132 4515 76188
rect 4515 76132 4519 76188
rect 4455 76128 4519 76132
rect 7479 76188 7543 76192
rect 7479 76132 7483 76188
rect 7483 76132 7539 76188
rect 7539 76132 7543 76188
rect 7479 76128 7543 76132
rect 7559 76188 7623 76192
rect 7559 76132 7563 76188
rect 7563 76132 7619 76188
rect 7619 76132 7623 76188
rect 7559 76128 7623 76132
rect 7639 76188 7703 76192
rect 7639 76132 7643 76188
rect 7643 76132 7699 76188
rect 7699 76132 7703 76188
rect 7639 76128 7703 76132
rect 7719 76188 7783 76192
rect 7719 76132 7723 76188
rect 7723 76132 7779 76188
rect 7779 76132 7783 76188
rect 7719 76128 7783 76132
rect 2584 75644 2648 75648
rect 2584 75588 2588 75644
rect 2588 75588 2644 75644
rect 2644 75588 2648 75644
rect 2584 75584 2648 75588
rect 2664 75644 2728 75648
rect 2664 75588 2668 75644
rect 2668 75588 2724 75644
rect 2724 75588 2728 75644
rect 2664 75584 2728 75588
rect 2744 75644 2808 75648
rect 2744 75588 2748 75644
rect 2748 75588 2804 75644
rect 2804 75588 2808 75644
rect 2744 75584 2808 75588
rect 2824 75644 2888 75648
rect 2824 75588 2828 75644
rect 2828 75588 2884 75644
rect 2884 75588 2888 75644
rect 2824 75584 2888 75588
rect 5847 75644 5911 75648
rect 5847 75588 5851 75644
rect 5851 75588 5907 75644
rect 5907 75588 5911 75644
rect 5847 75584 5911 75588
rect 5927 75644 5991 75648
rect 5927 75588 5931 75644
rect 5931 75588 5987 75644
rect 5987 75588 5991 75644
rect 5927 75584 5991 75588
rect 6007 75644 6071 75648
rect 6007 75588 6011 75644
rect 6011 75588 6067 75644
rect 6067 75588 6071 75644
rect 6007 75584 6071 75588
rect 6087 75644 6151 75648
rect 6087 75588 6091 75644
rect 6091 75588 6147 75644
rect 6147 75588 6151 75644
rect 6087 75584 6151 75588
rect 9111 75644 9175 75648
rect 9111 75588 9115 75644
rect 9115 75588 9171 75644
rect 9171 75588 9175 75644
rect 9111 75584 9175 75588
rect 9191 75644 9255 75648
rect 9191 75588 9195 75644
rect 9195 75588 9251 75644
rect 9251 75588 9255 75644
rect 9191 75584 9255 75588
rect 9271 75644 9335 75648
rect 9271 75588 9275 75644
rect 9275 75588 9331 75644
rect 9331 75588 9335 75644
rect 9271 75584 9335 75588
rect 9351 75644 9415 75648
rect 9351 75588 9355 75644
rect 9355 75588 9411 75644
rect 9411 75588 9415 75644
rect 9351 75584 9415 75588
rect 4215 75100 4279 75104
rect 4215 75044 4219 75100
rect 4219 75044 4275 75100
rect 4275 75044 4279 75100
rect 4215 75040 4279 75044
rect 4295 75100 4359 75104
rect 4295 75044 4299 75100
rect 4299 75044 4355 75100
rect 4355 75044 4359 75100
rect 4295 75040 4359 75044
rect 4375 75100 4439 75104
rect 4375 75044 4379 75100
rect 4379 75044 4435 75100
rect 4435 75044 4439 75100
rect 4375 75040 4439 75044
rect 4455 75100 4519 75104
rect 4455 75044 4459 75100
rect 4459 75044 4515 75100
rect 4515 75044 4519 75100
rect 4455 75040 4519 75044
rect 7479 75100 7543 75104
rect 7479 75044 7483 75100
rect 7483 75044 7539 75100
rect 7539 75044 7543 75100
rect 7479 75040 7543 75044
rect 7559 75100 7623 75104
rect 7559 75044 7563 75100
rect 7563 75044 7619 75100
rect 7619 75044 7623 75100
rect 7559 75040 7623 75044
rect 7639 75100 7703 75104
rect 7639 75044 7643 75100
rect 7643 75044 7699 75100
rect 7699 75044 7703 75100
rect 7639 75040 7703 75044
rect 7719 75100 7783 75104
rect 7719 75044 7723 75100
rect 7723 75044 7779 75100
rect 7779 75044 7783 75100
rect 7719 75040 7783 75044
rect 2584 74556 2648 74560
rect 2584 74500 2588 74556
rect 2588 74500 2644 74556
rect 2644 74500 2648 74556
rect 2584 74496 2648 74500
rect 2664 74556 2728 74560
rect 2664 74500 2668 74556
rect 2668 74500 2724 74556
rect 2724 74500 2728 74556
rect 2664 74496 2728 74500
rect 2744 74556 2808 74560
rect 2744 74500 2748 74556
rect 2748 74500 2804 74556
rect 2804 74500 2808 74556
rect 2744 74496 2808 74500
rect 2824 74556 2888 74560
rect 2824 74500 2828 74556
rect 2828 74500 2884 74556
rect 2884 74500 2888 74556
rect 2824 74496 2888 74500
rect 5847 74556 5911 74560
rect 5847 74500 5851 74556
rect 5851 74500 5907 74556
rect 5907 74500 5911 74556
rect 5847 74496 5911 74500
rect 5927 74556 5991 74560
rect 5927 74500 5931 74556
rect 5931 74500 5987 74556
rect 5987 74500 5991 74556
rect 5927 74496 5991 74500
rect 6007 74556 6071 74560
rect 6007 74500 6011 74556
rect 6011 74500 6067 74556
rect 6067 74500 6071 74556
rect 6007 74496 6071 74500
rect 6087 74556 6151 74560
rect 6087 74500 6091 74556
rect 6091 74500 6147 74556
rect 6147 74500 6151 74556
rect 6087 74496 6151 74500
rect 9111 74556 9175 74560
rect 9111 74500 9115 74556
rect 9115 74500 9171 74556
rect 9171 74500 9175 74556
rect 9111 74496 9175 74500
rect 9191 74556 9255 74560
rect 9191 74500 9195 74556
rect 9195 74500 9251 74556
rect 9251 74500 9255 74556
rect 9191 74496 9255 74500
rect 9271 74556 9335 74560
rect 9271 74500 9275 74556
rect 9275 74500 9331 74556
rect 9331 74500 9335 74556
rect 9271 74496 9335 74500
rect 9351 74556 9415 74560
rect 9351 74500 9355 74556
rect 9355 74500 9411 74556
rect 9411 74500 9415 74556
rect 9351 74496 9415 74500
rect 4215 74012 4279 74016
rect 4215 73956 4219 74012
rect 4219 73956 4275 74012
rect 4275 73956 4279 74012
rect 4215 73952 4279 73956
rect 4295 74012 4359 74016
rect 4295 73956 4299 74012
rect 4299 73956 4355 74012
rect 4355 73956 4359 74012
rect 4295 73952 4359 73956
rect 4375 74012 4439 74016
rect 4375 73956 4379 74012
rect 4379 73956 4435 74012
rect 4435 73956 4439 74012
rect 4375 73952 4439 73956
rect 4455 74012 4519 74016
rect 4455 73956 4459 74012
rect 4459 73956 4515 74012
rect 4515 73956 4519 74012
rect 4455 73952 4519 73956
rect 7479 74012 7543 74016
rect 7479 73956 7483 74012
rect 7483 73956 7539 74012
rect 7539 73956 7543 74012
rect 7479 73952 7543 73956
rect 7559 74012 7623 74016
rect 7559 73956 7563 74012
rect 7563 73956 7619 74012
rect 7619 73956 7623 74012
rect 7559 73952 7623 73956
rect 7639 74012 7703 74016
rect 7639 73956 7643 74012
rect 7643 73956 7699 74012
rect 7699 73956 7703 74012
rect 7639 73952 7703 73956
rect 7719 74012 7783 74016
rect 7719 73956 7723 74012
rect 7723 73956 7779 74012
rect 7779 73956 7783 74012
rect 7719 73952 7783 73956
rect 2584 73468 2648 73472
rect 2584 73412 2588 73468
rect 2588 73412 2644 73468
rect 2644 73412 2648 73468
rect 2584 73408 2648 73412
rect 2664 73468 2728 73472
rect 2664 73412 2668 73468
rect 2668 73412 2724 73468
rect 2724 73412 2728 73468
rect 2664 73408 2728 73412
rect 2744 73468 2808 73472
rect 2744 73412 2748 73468
rect 2748 73412 2804 73468
rect 2804 73412 2808 73468
rect 2744 73408 2808 73412
rect 2824 73468 2888 73472
rect 2824 73412 2828 73468
rect 2828 73412 2884 73468
rect 2884 73412 2888 73468
rect 2824 73408 2888 73412
rect 5847 73468 5911 73472
rect 5847 73412 5851 73468
rect 5851 73412 5907 73468
rect 5907 73412 5911 73468
rect 5847 73408 5911 73412
rect 5927 73468 5991 73472
rect 5927 73412 5931 73468
rect 5931 73412 5987 73468
rect 5987 73412 5991 73468
rect 5927 73408 5991 73412
rect 6007 73468 6071 73472
rect 6007 73412 6011 73468
rect 6011 73412 6067 73468
rect 6067 73412 6071 73468
rect 6007 73408 6071 73412
rect 6087 73468 6151 73472
rect 6087 73412 6091 73468
rect 6091 73412 6147 73468
rect 6147 73412 6151 73468
rect 6087 73408 6151 73412
rect 9111 73468 9175 73472
rect 9111 73412 9115 73468
rect 9115 73412 9171 73468
rect 9171 73412 9175 73468
rect 9111 73408 9175 73412
rect 9191 73468 9255 73472
rect 9191 73412 9195 73468
rect 9195 73412 9251 73468
rect 9251 73412 9255 73468
rect 9191 73408 9255 73412
rect 9271 73468 9335 73472
rect 9271 73412 9275 73468
rect 9275 73412 9331 73468
rect 9331 73412 9335 73468
rect 9271 73408 9335 73412
rect 9351 73468 9415 73472
rect 9351 73412 9355 73468
rect 9355 73412 9411 73468
rect 9411 73412 9415 73468
rect 9351 73408 9415 73412
rect 4215 72924 4279 72928
rect 4215 72868 4219 72924
rect 4219 72868 4275 72924
rect 4275 72868 4279 72924
rect 4215 72864 4279 72868
rect 4295 72924 4359 72928
rect 4295 72868 4299 72924
rect 4299 72868 4355 72924
rect 4355 72868 4359 72924
rect 4295 72864 4359 72868
rect 4375 72924 4439 72928
rect 4375 72868 4379 72924
rect 4379 72868 4435 72924
rect 4435 72868 4439 72924
rect 4375 72864 4439 72868
rect 4455 72924 4519 72928
rect 4455 72868 4459 72924
rect 4459 72868 4515 72924
rect 4515 72868 4519 72924
rect 4455 72864 4519 72868
rect 7479 72924 7543 72928
rect 7479 72868 7483 72924
rect 7483 72868 7539 72924
rect 7539 72868 7543 72924
rect 7479 72864 7543 72868
rect 7559 72924 7623 72928
rect 7559 72868 7563 72924
rect 7563 72868 7619 72924
rect 7619 72868 7623 72924
rect 7559 72864 7623 72868
rect 7639 72924 7703 72928
rect 7639 72868 7643 72924
rect 7643 72868 7699 72924
rect 7699 72868 7703 72924
rect 7639 72864 7703 72868
rect 7719 72924 7783 72928
rect 7719 72868 7723 72924
rect 7723 72868 7779 72924
rect 7779 72868 7783 72924
rect 7719 72864 7783 72868
rect 2584 72380 2648 72384
rect 2584 72324 2588 72380
rect 2588 72324 2644 72380
rect 2644 72324 2648 72380
rect 2584 72320 2648 72324
rect 2664 72380 2728 72384
rect 2664 72324 2668 72380
rect 2668 72324 2724 72380
rect 2724 72324 2728 72380
rect 2664 72320 2728 72324
rect 2744 72380 2808 72384
rect 2744 72324 2748 72380
rect 2748 72324 2804 72380
rect 2804 72324 2808 72380
rect 2744 72320 2808 72324
rect 2824 72380 2888 72384
rect 2824 72324 2828 72380
rect 2828 72324 2884 72380
rect 2884 72324 2888 72380
rect 2824 72320 2888 72324
rect 5847 72380 5911 72384
rect 5847 72324 5851 72380
rect 5851 72324 5907 72380
rect 5907 72324 5911 72380
rect 5847 72320 5911 72324
rect 5927 72380 5991 72384
rect 5927 72324 5931 72380
rect 5931 72324 5987 72380
rect 5987 72324 5991 72380
rect 5927 72320 5991 72324
rect 6007 72380 6071 72384
rect 6007 72324 6011 72380
rect 6011 72324 6067 72380
rect 6067 72324 6071 72380
rect 6007 72320 6071 72324
rect 6087 72380 6151 72384
rect 6087 72324 6091 72380
rect 6091 72324 6147 72380
rect 6147 72324 6151 72380
rect 6087 72320 6151 72324
rect 9111 72380 9175 72384
rect 9111 72324 9115 72380
rect 9115 72324 9171 72380
rect 9171 72324 9175 72380
rect 9111 72320 9175 72324
rect 9191 72380 9255 72384
rect 9191 72324 9195 72380
rect 9195 72324 9251 72380
rect 9251 72324 9255 72380
rect 9191 72320 9255 72324
rect 9271 72380 9335 72384
rect 9271 72324 9275 72380
rect 9275 72324 9331 72380
rect 9331 72324 9335 72380
rect 9271 72320 9335 72324
rect 9351 72380 9415 72384
rect 9351 72324 9355 72380
rect 9355 72324 9411 72380
rect 9411 72324 9415 72380
rect 9351 72320 9415 72324
rect 4215 71836 4279 71840
rect 4215 71780 4219 71836
rect 4219 71780 4275 71836
rect 4275 71780 4279 71836
rect 4215 71776 4279 71780
rect 4295 71836 4359 71840
rect 4295 71780 4299 71836
rect 4299 71780 4355 71836
rect 4355 71780 4359 71836
rect 4295 71776 4359 71780
rect 4375 71836 4439 71840
rect 4375 71780 4379 71836
rect 4379 71780 4435 71836
rect 4435 71780 4439 71836
rect 4375 71776 4439 71780
rect 4455 71836 4519 71840
rect 4455 71780 4459 71836
rect 4459 71780 4515 71836
rect 4515 71780 4519 71836
rect 4455 71776 4519 71780
rect 7479 71836 7543 71840
rect 7479 71780 7483 71836
rect 7483 71780 7539 71836
rect 7539 71780 7543 71836
rect 7479 71776 7543 71780
rect 7559 71836 7623 71840
rect 7559 71780 7563 71836
rect 7563 71780 7619 71836
rect 7619 71780 7623 71836
rect 7559 71776 7623 71780
rect 7639 71836 7703 71840
rect 7639 71780 7643 71836
rect 7643 71780 7699 71836
rect 7699 71780 7703 71836
rect 7639 71776 7703 71780
rect 7719 71836 7783 71840
rect 7719 71780 7723 71836
rect 7723 71780 7779 71836
rect 7779 71780 7783 71836
rect 7719 71776 7783 71780
rect 2584 71292 2648 71296
rect 2584 71236 2588 71292
rect 2588 71236 2644 71292
rect 2644 71236 2648 71292
rect 2584 71232 2648 71236
rect 2664 71292 2728 71296
rect 2664 71236 2668 71292
rect 2668 71236 2724 71292
rect 2724 71236 2728 71292
rect 2664 71232 2728 71236
rect 2744 71292 2808 71296
rect 2744 71236 2748 71292
rect 2748 71236 2804 71292
rect 2804 71236 2808 71292
rect 2744 71232 2808 71236
rect 2824 71292 2888 71296
rect 2824 71236 2828 71292
rect 2828 71236 2884 71292
rect 2884 71236 2888 71292
rect 2824 71232 2888 71236
rect 5847 71292 5911 71296
rect 5847 71236 5851 71292
rect 5851 71236 5907 71292
rect 5907 71236 5911 71292
rect 5847 71232 5911 71236
rect 5927 71292 5991 71296
rect 5927 71236 5931 71292
rect 5931 71236 5987 71292
rect 5987 71236 5991 71292
rect 5927 71232 5991 71236
rect 6007 71292 6071 71296
rect 6007 71236 6011 71292
rect 6011 71236 6067 71292
rect 6067 71236 6071 71292
rect 6007 71232 6071 71236
rect 6087 71292 6151 71296
rect 6087 71236 6091 71292
rect 6091 71236 6147 71292
rect 6147 71236 6151 71292
rect 6087 71232 6151 71236
rect 9111 71292 9175 71296
rect 9111 71236 9115 71292
rect 9115 71236 9171 71292
rect 9171 71236 9175 71292
rect 9111 71232 9175 71236
rect 9191 71292 9255 71296
rect 9191 71236 9195 71292
rect 9195 71236 9251 71292
rect 9251 71236 9255 71292
rect 9191 71232 9255 71236
rect 9271 71292 9335 71296
rect 9271 71236 9275 71292
rect 9275 71236 9331 71292
rect 9331 71236 9335 71292
rect 9271 71232 9335 71236
rect 9351 71292 9415 71296
rect 9351 71236 9355 71292
rect 9355 71236 9411 71292
rect 9411 71236 9415 71292
rect 9351 71232 9415 71236
rect 4215 70748 4279 70752
rect 4215 70692 4219 70748
rect 4219 70692 4275 70748
rect 4275 70692 4279 70748
rect 4215 70688 4279 70692
rect 4295 70748 4359 70752
rect 4295 70692 4299 70748
rect 4299 70692 4355 70748
rect 4355 70692 4359 70748
rect 4295 70688 4359 70692
rect 4375 70748 4439 70752
rect 4375 70692 4379 70748
rect 4379 70692 4435 70748
rect 4435 70692 4439 70748
rect 4375 70688 4439 70692
rect 4455 70748 4519 70752
rect 4455 70692 4459 70748
rect 4459 70692 4515 70748
rect 4515 70692 4519 70748
rect 4455 70688 4519 70692
rect 7479 70748 7543 70752
rect 7479 70692 7483 70748
rect 7483 70692 7539 70748
rect 7539 70692 7543 70748
rect 7479 70688 7543 70692
rect 7559 70748 7623 70752
rect 7559 70692 7563 70748
rect 7563 70692 7619 70748
rect 7619 70692 7623 70748
rect 7559 70688 7623 70692
rect 7639 70748 7703 70752
rect 7639 70692 7643 70748
rect 7643 70692 7699 70748
rect 7699 70692 7703 70748
rect 7639 70688 7703 70692
rect 7719 70748 7783 70752
rect 7719 70692 7723 70748
rect 7723 70692 7779 70748
rect 7779 70692 7783 70748
rect 7719 70688 7783 70692
rect 2584 70204 2648 70208
rect 2584 70148 2588 70204
rect 2588 70148 2644 70204
rect 2644 70148 2648 70204
rect 2584 70144 2648 70148
rect 2664 70204 2728 70208
rect 2664 70148 2668 70204
rect 2668 70148 2724 70204
rect 2724 70148 2728 70204
rect 2664 70144 2728 70148
rect 2744 70204 2808 70208
rect 2744 70148 2748 70204
rect 2748 70148 2804 70204
rect 2804 70148 2808 70204
rect 2744 70144 2808 70148
rect 2824 70204 2888 70208
rect 2824 70148 2828 70204
rect 2828 70148 2884 70204
rect 2884 70148 2888 70204
rect 2824 70144 2888 70148
rect 5847 70204 5911 70208
rect 5847 70148 5851 70204
rect 5851 70148 5907 70204
rect 5907 70148 5911 70204
rect 5847 70144 5911 70148
rect 5927 70204 5991 70208
rect 5927 70148 5931 70204
rect 5931 70148 5987 70204
rect 5987 70148 5991 70204
rect 5927 70144 5991 70148
rect 6007 70204 6071 70208
rect 6007 70148 6011 70204
rect 6011 70148 6067 70204
rect 6067 70148 6071 70204
rect 6007 70144 6071 70148
rect 6087 70204 6151 70208
rect 6087 70148 6091 70204
rect 6091 70148 6147 70204
rect 6147 70148 6151 70204
rect 6087 70144 6151 70148
rect 9111 70204 9175 70208
rect 9111 70148 9115 70204
rect 9115 70148 9171 70204
rect 9171 70148 9175 70204
rect 9111 70144 9175 70148
rect 9191 70204 9255 70208
rect 9191 70148 9195 70204
rect 9195 70148 9251 70204
rect 9251 70148 9255 70204
rect 9191 70144 9255 70148
rect 9271 70204 9335 70208
rect 9271 70148 9275 70204
rect 9275 70148 9331 70204
rect 9331 70148 9335 70204
rect 9271 70144 9335 70148
rect 9351 70204 9415 70208
rect 9351 70148 9355 70204
rect 9355 70148 9411 70204
rect 9411 70148 9415 70204
rect 9351 70144 9415 70148
rect 4215 69660 4279 69664
rect 4215 69604 4219 69660
rect 4219 69604 4275 69660
rect 4275 69604 4279 69660
rect 4215 69600 4279 69604
rect 4295 69660 4359 69664
rect 4295 69604 4299 69660
rect 4299 69604 4355 69660
rect 4355 69604 4359 69660
rect 4295 69600 4359 69604
rect 4375 69660 4439 69664
rect 4375 69604 4379 69660
rect 4379 69604 4435 69660
rect 4435 69604 4439 69660
rect 4375 69600 4439 69604
rect 4455 69660 4519 69664
rect 4455 69604 4459 69660
rect 4459 69604 4515 69660
rect 4515 69604 4519 69660
rect 4455 69600 4519 69604
rect 7479 69660 7543 69664
rect 7479 69604 7483 69660
rect 7483 69604 7539 69660
rect 7539 69604 7543 69660
rect 7479 69600 7543 69604
rect 7559 69660 7623 69664
rect 7559 69604 7563 69660
rect 7563 69604 7619 69660
rect 7619 69604 7623 69660
rect 7559 69600 7623 69604
rect 7639 69660 7703 69664
rect 7639 69604 7643 69660
rect 7643 69604 7699 69660
rect 7699 69604 7703 69660
rect 7639 69600 7703 69604
rect 7719 69660 7783 69664
rect 7719 69604 7723 69660
rect 7723 69604 7779 69660
rect 7779 69604 7783 69660
rect 7719 69600 7783 69604
rect 2584 69116 2648 69120
rect 2584 69060 2588 69116
rect 2588 69060 2644 69116
rect 2644 69060 2648 69116
rect 2584 69056 2648 69060
rect 2664 69116 2728 69120
rect 2664 69060 2668 69116
rect 2668 69060 2724 69116
rect 2724 69060 2728 69116
rect 2664 69056 2728 69060
rect 2744 69116 2808 69120
rect 2744 69060 2748 69116
rect 2748 69060 2804 69116
rect 2804 69060 2808 69116
rect 2744 69056 2808 69060
rect 2824 69116 2888 69120
rect 2824 69060 2828 69116
rect 2828 69060 2884 69116
rect 2884 69060 2888 69116
rect 2824 69056 2888 69060
rect 5847 69116 5911 69120
rect 5847 69060 5851 69116
rect 5851 69060 5907 69116
rect 5907 69060 5911 69116
rect 5847 69056 5911 69060
rect 5927 69116 5991 69120
rect 5927 69060 5931 69116
rect 5931 69060 5987 69116
rect 5987 69060 5991 69116
rect 5927 69056 5991 69060
rect 6007 69116 6071 69120
rect 6007 69060 6011 69116
rect 6011 69060 6067 69116
rect 6067 69060 6071 69116
rect 6007 69056 6071 69060
rect 6087 69116 6151 69120
rect 6087 69060 6091 69116
rect 6091 69060 6147 69116
rect 6147 69060 6151 69116
rect 6087 69056 6151 69060
rect 9111 69116 9175 69120
rect 9111 69060 9115 69116
rect 9115 69060 9171 69116
rect 9171 69060 9175 69116
rect 9111 69056 9175 69060
rect 9191 69116 9255 69120
rect 9191 69060 9195 69116
rect 9195 69060 9251 69116
rect 9251 69060 9255 69116
rect 9191 69056 9255 69060
rect 9271 69116 9335 69120
rect 9271 69060 9275 69116
rect 9275 69060 9331 69116
rect 9331 69060 9335 69116
rect 9271 69056 9335 69060
rect 9351 69116 9415 69120
rect 9351 69060 9355 69116
rect 9355 69060 9411 69116
rect 9411 69060 9415 69116
rect 9351 69056 9415 69060
rect 1164 68988 1228 69052
rect 4215 68572 4279 68576
rect 4215 68516 4219 68572
rect 4219 68516 4275 68572
rect 4275 68516 4279 68572
rect 4215 68512 4279 68516
rect 4295 68572 4359 68576
rect 4295 68516 4299 68572
rect 4299 68516 4355 68572
rect 4355 68516 4359 68572
rect 4295 68512 4359 68516
rect 4375 68572 4439 68576
rect 4375 68516 4379 68572
rect 4379 68516 4435 68572
rect 4435 68516 4439 68572
rect 4375 68512 4439 68516
rect 4455 68572 4519 68576
rect 4455 68516 4459 68572
rect 4459 68516 4515 68572
rect 4515 68516 4519 68572
rect 4455 68512 4519 68516
rect 7479 68572 7543 68576
rect 7479 68516 7483 68572
rect 7483 68516 7539 68572
rect 7539 68516 7543 68572
rect 7479 68512 7543 68516
rect 7559 68572 7623 68576
rect 7559 68516 7563 68572
rect 7563 68516 7619 68572
rect 7619 68516 7623 68572
rect 7559 68512 7623 68516
rect 7639 68572 7703 68576
rect 7639 68516 7643 68572
rect 7643 68516 7699 68572
rect 7699 68516 7703 68572
rect 7639 68512 7703 68516
rect 7719 68572 7783 68576
rect 7719 68516 7723 68572
rect 7723 68516 7779 68572
rect 7779 68516 7783 68572
rect 7719 68512 7783 68516
rect 2584 68028 2648 68032
rect 2584 67972 2588 68028
rect 2588 67972 2644 68028
rect 2644 67972 2648 68028
rect 2584 67968 2648 67972
rect 2664 68028 2728 68032
rect 2664 67972 2668 68028
rect 2668 67972 2724 68028
rect 2724 67972 2728 68028
rect 2664 67968 2728 67972
rect 2744 68028 2808 68032
rect 2744 67972 2748 68028
rect 2748 67972 2804 68028
rect 2804 67972 2808 68028
rect 2744 67968 2808 67972
rect 2824 68028 2888 68032
rect 2824 67972 2828 68028
rect 2828 67972 2884 68028
rect 2884 67972 2888 68028
rect 2824 67968 2888 67972
rect 5847 68028 5911 68032
rect 5847 67972 5851 68028
rect 5851 67972 5907 68028
rect 5907 67972 5911 68028
rect 5847 67968 5911 67972
rect 5927 68028 5991 68032
rect 5927 67972 5931 68028
rect 5931 67972 5987 68028
rect 5987 67972 5991 68028
rect 5927 67968 5991 67972
rect 6007 68028 6071 68032
rect 6007 67972 6011 68028
rect 6011 67972 6067 68028
rect 6067 67972 6071 68028
rect 6007 67968 6071 67972
rect 6087 68028 6151 68032
rect 6087 67972 6091 68028
rect 6091 67972 6147 68028
rect 6147 67972 6151 68028
rect 6087 67968 6151 67972
rect 9111 68028 9175 68032
rect 9111 67972 9115 68028
rect 9115 67972 9171 68028
rect 9171 67972 9175 68028
rect 9111 67968 9175 67972
rect 9191 68028 9255 68032
rect 9191 67972 9195 68028
rect 9195 67972 9251 68028
rect 9251 67972 9255 68028
rect 9191 67968 9255 67972
rect 9271 68028 9335 68032
rect 9271 67972 9275 68028
rect 9275 67972 9331 68028
rect 9331 67972 9335 68028
rect 9271 67968 9335 67972
rect 9351 68028 9415 68032
rect 9351 67972 9355 68028
rect 9355 67972 9411 68028
rect 9411 67972 9415 68028
rect 9351 67968 9415 67972
rect 4215 67484 4279 67488
rect 4215 67428 4219 67484
rect 4219 67428 4275 67484
rect 4275 67428 4279 67484
rect 4215 67424 4279 67428
rect 4295 67484 4359 67488
rect 4295 67428 4299 67484
rect 4299 67428 4355 67484
rect 4355 67428 4359 67484
rect 4295 67424 4359 67428
rect 4375 67484 4439 67488
rect 4375 67428 4379 67484
rect 4379 67428 4435 67484
rect 4435 67428 4439 67484
rect 4375 67424 4439 67428
rect 4455 67484 4519 67488
rect 4455 67428 4459 67484
rect 4459 67428 4515 67484
rect 4515 67428 4519 67484
rect 4455 67424 4519 67428
rect 7479 67484 7543 67488
rect 7479 67428 7483 67484
rect 7483 67428 7539 67484
rect 7539 67428 7543 67484
rect 7479 67424 7543 67428
rect 7559 67484 7623 67488
rect 7559 67428 7563 67484
rect 7563 67428 7619 67484
rect 7619 67428 7623 67484
rect 7559 67424 7623 67428
rect 7639 67484 7703 67488
rect 7639 67428 7643 67484
rect 7643 67428 7699 67484
rect 7699 67428 7703 67484
rect 7639 67424 7703 67428
rect 7719 67484 7783 67488
rect 7719 67428 7723 67484
rect 7723 67428 7779 67484
rect 7779 67428 7783 67484
rect 7719 67424 7783 67428
rect 2584 66940 2648 66944
rect 2584 66884 2588 66940
rect 2588 66884 2644 66940
rect 2644 66884 2648 66940
rect 2584 66880 2648 66884
rect 2664 66940 2728 66944
rect 2664 66884 2668 66940
rect 2668 66884 2724 66940
rect 2724 66884 2728 66940
rect 2664 66880 2728 66884
rect 2744 66940 2808 66944
rect 2744 66884 2748 66940
rect 2748 66884 2804 66940
rect 2804 66884 2808 66940
rect 2744 66880 2808 66884
rect 2824 66940 2888 66944
rect 2824 66884 2828 66940
rect 2828 66884 2884 66940
rect 2884 66884 2888 66940
rect 2824 66880 2888 66884
rect 5847 66940 5911 66944
rect 5847 66884 5851 66940
rect 5851 66884 5907 66940
rect 5907 66884 5911 66940
rect 5847 66880 5911 66884
rect 5927 66940 5991 66944
rect 5927 66884 5931 66940
rect 5931 66884 5987 66940
rect 5987 66884 5991 66940
rect 5927 66880 5991 66884
rect 6007 66940 6071 66944
rect 6007 66884 6011 66940
rect 6011 66884 6067 66940
rect 6067 66884 6071 66940
rect 6007 66880 6071 66884
rect 6087 66940 6151 66944
rect 6087 66884 6091 66940
rect 6091 66884 6147 66940
rect 6147 66884 6151 66940
rect 6087 66880 6151 66884
rect 9111 66940 9175 66944
rect 9111 66884 9115 66940
rect 9115 66884 9171 66940
rect 9171 66884 9175 66940
rect 9111 66880 9175 66884
rect 9191 66940 9255 66944
rect 9191 66884 9195 66940
rect 9195 66884 9251 66940
rect 9251 66884 9255 66940
rect 9191 66880 9255 66884
rect 9271 66940 9335 66944
rect 9271 66884 9275 66940
rect 9275 66884 9331 66940
rect 9331 66884 9335 66940
rect 9271 66880 9335 66884
rect 9351 66940 9415 66944
rect 9351 66884 9355 66940
rect 9355 66884 9411 66940
rect 9411 66884 9415 66940
rect 9351 66880 9415 66884
rect 4215 66396 4279 66400
rect 4215 66340 4219 66396
rect 4219 66340 4275 66396
rect 4275 66340 4279 66396
rect 4215 66336 4279 66340
rect 4295 66396 4359 66400
rect 4295 66340 4299 66396
rect 4299 66340 4355 66396
rect 4355 66340 4359 66396
rect 4295 66336 4359 66340
rect 4375 66396 4439 66400
rect 4375 66340 4379 66396
rect 4379 66340 4435 66396
rect 4435 66340 4439 66396
rect 4375 66336 4439 66340
rect 4455 66396 4519 66400
rect 4455 66340 4459 66396
rect 4459 66340 4515 66396
rect 4515 66340 4519 66396
rect 4455 66336 4519 66340
rect 7479 66396 7543 66400
rect 7479 66340 7483 66396
rect 7483 66340 7539 66396
rect 7539 66340 7543 66396
rect 7479 66336 7543 66340
rect 7559 66396 7623 66400
rect 7559 66340 7563 66396
rect 7563 66340 7619 66396
rect 7619 66340 7623 66396
rect 7559 66336 7623 66340
rect 7639 66396 7703 66400
rect 7639 66340 7643 66396
rect 7643 66340 7699 66396
rect 7699 66340 7703 66396
rect 7639 66336 7703 66340
rect 7719 66396 7783 66400
rect 7719 66340 7723 66396
rect 7723 66340 7779 66396
rect 7779 66340 7783 66396
rect 7719 66336 7783 66340
rect 2584 65852 2648 65856
rect 2584 65796 2588 65852
rect 2588 65796 2644 65852
rect 2644 65796 2648 65852
rect 2584 65792 2648 65796
rect 2664 65852 2728 65856
rect 2664 65796 2668 65852
rect 2668 65796 2724 65852
rect 2724 65796 2728 65852
rect 2664 65792 2728 65796
rect 2744 65852 2808 65856
rect 2744 65796 2748 65852
rect 2748 65796 2804 65852
rect 2804 65796 2808 65852
rect 2744 65792 2808 65796
rect 2824 65852 2888 65856
rect 2824 65796 2828 65852
rect 2828 65796 2884 65852
rect 2884 65796 2888 65852
rect 2824 65792 2888 65796
rect 5847 65852 5911 65856
rect 5847 65796 5851 65852
rect 5851 65796 5907 65852
rect 5907 65796 5911 65852
rect 5847 65792 5911 65796
rect 5927 65852 5991 65856
rect 5927 65796 5931 65852
rect 5931 65796 5987 65852
rect 5987 65796 5991 65852
rect 5927 65792 5991 65796
rect 6007 65852 6071 65856
rect 6007 65796 6011 65852
rect 6011 65796 6067 65852
rect 6067 65796 6071 65852
rect 6007 65792 6071 65796
rect 6087 65852 6151 65856
rect 6087 65796 6091 65852
rect 6091 65796 6147 65852
rect 6147 65796 6151 65852
rect 6087 65792 6151 65796
rect 9111 65852 9175 65856
rect 9111 65796 9115 65852
rect 9115 65796 9171 65852
rect 9171 65796 9175 65852
rect 9111 65792 9175 65796
rect 9191 65852 9255 65856
rect 9191 65796 9195 65852
rect 9195 65796 9251 65852
rect 9251 65796 9255 65852
rect 9191 65792 9255 65796
rect 9271 65852 9335 65856
rect 9271 65796 9275 65852
rect 9275 65796 9331 65852
rect 9331 65796 9335 65852
rect 9271 65792 9335 65796
rect 9351 65852 9415 65856
rect 9351 65796 9355 65852
rect 9355 65796 9411 65852
rect 9411 65796 9415 65852
rect 9351 65792 9415 65796
rect 4215 65308 4279 65312
rect 4215 65252 4219 65308
rect 4219 65252 4275 65308
rect 4275 65252 4279 65308
rect 4215 65248 4279 65252
rect 4295 65308 4359 65312
rect 4295 65252 4299 65308
rect 4299 65252 4355 65308
rect 4355 65252 4359 65308
rect 4295 65248 4359 65252
rect 4375 65308 4439 65312
rect 4375 65252 4379 65308
rect 4379 65252 4435 65308
rect 4435 65252 4439 65308
rect 4375 65248 4439 65252
rect 4455 65308 4519 65312
rect 4455 65252 4459 65308
rect 4459 65252 4515 65308
rect 4515 65252 4519 65308
rect 4455 65248 4519 65252
rect 7479 65308 7543 65312
rect 7479 65252 7483 65308
rect 7483 65252 7539 65308
rect 7539 65252 7543 65308
rect 7479 65248 7543 65252
rect 7559 65308 7623 65312
rect 7559 65252 7563 65308
rect 7563 65252 7619 65308
rect 7619 65252 7623 65308
rect 7559 65248 7623 65252
rect 7639 65308 7703 65312
rect 7639 65252 7643 65308
rect 7643 65252 7699 65308
rect 7699 65252 7703 65308
rect 7639 65248 7703 65252
rect 7719 65308 7783 65312
rect 7719 65252 7723 65308
rect 7723 65252 7779 65308
rect 7779 65252 7783 65308
rect 7719 65248 7783 65252
rect 2584 64764 2648 64768
rect 2584 64708 2588 64764
rect 2588 64708 2644 64764
rect 2644 64708 2648 64764
rect 2584 64704 2648 64708
rect 2664 64764 2728 64768
rect 2664 64708 2668 64764
rect 2668 64708 2724 64764
rect 2724 64708 2728 64764
rect 2664 64704 2728 64708
rect 2744 64764 2808 64768
rect 2744 64708 2748 64764
rect 2748 64708 2804 64764
rect 2804 64708 2808 64764
rect 2744 64704 2808 64708
rect 2824 64764 2888 64768
rect 2824 64708 2828 64764
rect 2828 64708 2884 64764
rect 2884 64708 2888 64764
rect 2824 64704 2888 64708
rect 5847 64764 5911 64768
rect 5847 64708 5851 64764
rect 5851 64708 5907 64764
rect 5907 64708 5911 64764
rect 5847 64704 5911 64708
rect 5927 64764 5991 64768
rect 5927 64708 5931 64764
rect 5931 64708 5987 64764
rect 5987 64708 5991 64764
rect 5927 64704 5991 64708
rect 6007 64764 6071 64768
rect 6007 64708 6011 64764
rect 6011 64708 6067 64764
rect 6067 64708 6071 64764
rect 6007 64704 6071 64708
rect 6087 64764 6151 64768
rect 6087 64708 6091 64764
rect 6091 64708 6147 64764
rect 6147 64708 6151 64764
rect 6087 64704 6151 64708
rect 9111 64764 9175 64768
rect 9111 64708 9115 64764
rect 9115 64708 9171 64764
rect 9171 64708 9175 64764
rect 9111 64704 9175 64708
rect 9191 64764 9255 64768
rect 9191 64708 9195 64764
rect 9195 64708 9251 64764
rect 9251 64708 9255 64764
rect 9191 64704 9255 64708
rect 9271 64764 9335 64768
rect 9271 64708 9275 64764
rect 9275 64708 9331 64764
rect 9331 64708 9335 64764
rect 9271 64704 9335 64708
rect 9351 64764 9415 64768
rect 9351 64708 9355 64764
rect 9355 64708 9411 64764
rect 9411 64708 9415 64764
rect 9351 64704 9415 64708
rect 4215 64220 4279 64224
rect 4215 64164 4219 64220
rect 4219 64164 4275 64220
rect 4275 64164 4279 64220
rect 4215 64160 4279 64164
rect 4295 64220 4359 64224
rect 4295 64164 4299 64220
rect 4299 64164 4355 64220
rect 4355 64164 4359 64220
rect 4295 64160 4359 64164
rect 4375 64220 4439 64224
rect 4375 64164 4379 64220
rect 4379 64164 4435 64220
rect 4435 64164 4439 64220
rect 4375 64160 4439 64164
rect 4455 64220 4519 64224
rect 4455 64164 4459 64220
rect 4459 64164 4515 64220
rect 4515 64164 4519 64220
rect 4455 64160 4519 64164
rect 7479 64220 7543 64224
rect 7479 64164 7483 64220
rect 7483 64164 7539 64220
rect 7539 64164 7543 64220
rect 7479 64160 7543 64164
rect 7559 64220 7623 64224
rect 7559 64164 7563 64220
rect 7563 64164 7619 64220
rect 7619 64164 7623 64220
rect 7559 64160 7623 64164
rect 7639 64220 7703 64224
rect 7639 64164 7643 64220
rect 7643 64164 7699 64220
rect 7699 64164 7703 64220
rect 7639 64160 7703 64164
rect 7719 64220 7783 64224
rect 7719 64164 7723 64220
rect 7723 64164 7779 64220
rect 7779 64164 7783 64220
rect 7719 64160 7783 64164
rect 2584 63676 2648 63680
rect 2584 63620 2588 63676
rect 2588 63620 2644 63676
rect 2644 63620 2648 63676
rect 2584 63616 2648 63620
rect 2664 63676 2728 63680
rect 2664 63620 2668 63676
rect 2668 63620 2724 63676
rect 2724 63620 2728 63676
rect 2664 63616 2728 63620
rect 2744 63676 2808 63680
rect 2744 63620 2748 63676
rect 2748 63620 2804 63676
rect 2804 63620 2808 63676
rect 2744 63616 2808 63620
rect 2824 63676 2888 63680
rect 2824 63620 2828 63676
rect 2828 63620 2884 63676
rect 2884 63620 2888 63676
rect 2824 63616 2888 63620
rect 5847 63676 5911 63680
rect 5847 63620 5851 63676
rect 5851 63620 5907 63676
rect 5907 63620 5911 63676
rect 5847 63616 5911 63620
rect 5927 63676 5991 63680
rect 5927 63620 5931 63676
rect 5931 63620 5987 63676
rect 5987 63620 5991 63676
rect 5927 63616 5991 63620
rect 6007 63676 6071 63680
rect 6007 63620 6011 63676
rect 6011 63620 6067 63676
rect 6067 63620 6071 63676
rect 6007 63616 6071 63620
rect 6087 63676 6151 63680
rect 6087 63620 6091 63676
rect 6091 63620 6147 63676
rect 6147 63620 6151 63676
rect 6087 63616 6151 63620
rect 9111 63676 9175 63680
rect 9111 63620 9115 63676
rect 9115 63620 9171 63676
rect 9171 63620 9175 63676
rect 9111 63616 9175 63620
rect 9191 63676 9255 63680
rect 9191 63620 9195 63676
rect 9195 63620 9251 63676
rect 9251 63620 9255 63676
rect 9191 63616 9255 63620
rect 9271 63676 9335 63680
rect 9271 63620 9275 63676
rect 9275 63620 9331 63676
rect 9331 63620 9335 63676
rect 9271 63616 9335 63620
rect 9351 63676 9415 63680
rect 9351 63620 9355 63676
rect 9355 63620 9411 63676
rect 9411 63620 9415 63676
rect 9351 63616 9415 63620
rect 4215 63132 4279 63136
rect 4215 63076 4219 63132
rect 4219 63076 4275 63132
rect 4275 63076 4279 63132
rect 4215 63072 4279 63076
rect 4295 63132 4359 63136
rect 4295 63076 4299 63132
rect 4299 63076 4355 63132
rect 4355 63076 4359 63132
rect 4295 63072 4359 63076
rect 4375 63132 4439 63136
rect 4375 63076 4379 63132
rect 4379 63076 4435 63132
rect 4435 63076 4439 63132
rect 4375 63072 4439 63076
rect 4455 63132 4519 63136
rect 4455 63076 4459 63132
rect 4459 63076 4515 63132
rect 4515 63076 4519 63132
rect 4455 63072 4519 63076
rect 7479 63132 7543 63136
rect 7479 63076 7483 63132
rect 7483 63076 7539 63132
rect 7539 63076 7543 63132
rect 7479 63072 7543 63076
rect 7559 63132 7623 63136
rect 7559 63076 7563 63132
rect 7563 63076 7619 63132
rect 7619 63076 7623 63132
rect 7559 63072 7623 63076
rect 7639 63132 7703 63136
rect 7639 63076 7643 63132
rect 7643 63076 7699 63132
rect 7699 63076 7703 63132
rect 7639 63072 7703 63076
rect 7719 63132 7783 63136
rect 7719 63076 7723 63132
rect 7723 63076 7779 63132
rect 7779 63076 7783 63132
rect 7719 63072 7783 63076
rect 2584 62588 2648 62592
rect 2584 62532 2588 62588
rect 2588 62532 2644 62588
rect 2644 62532 2648 62588
rect 2584 62528 2648 62532
rect 2664 62588 2728 62592
rect 2664 62532 2668 62588
rect 2668 62532 2724 62588
rect 2724 62532 2728 62588
rect 2664 62528 2728 62532
rect 2744 62588 2808 62592
rect 2744 62532 2748 62588
rect 2748 62532 2804 62588
rect 2804 62532 2808 62588
rect 2744 62528 2808 62532
rect 2824 62588 2888 62592
rect 2824 62532 2828 62588
rect 2828 62532 2884 62588
rect 2884 62532 2888 62588
rect 2824 62528 2888 62532
rect 5847 62588 5911 62592
rect 5847 62532 5851 62588
rect 5851 62532 5907 62588
rect 5907 62532 5911 62588
rect 5847 62528 5911 62532
rect 5927 62588 5991 62592
rect 5927 62532 5931 62588
rect 5931 62532 5987 62588
rect 5987 62532 5991 62588
rect 5927 62528 5991 62532
rect 6007 62588 6071 62592
rect 6007 62532 6011 62588
rect 6011 62532 6067 62588
rect 6067 62532 6071 62588
rect 6007 62528 6071 62532
rect 6087 62588 6151 62592
rect 6087 62532 6091 62588
rect 6091 62532 6147 62588
rect 6147 62532 6151 62588
rect 6087 62528 6151 62532
rect 9111 62588 9175 62592
rect 9111 62532 9115 62588
rect 9115 62532 9171 62588
rect 9171 62532 9175 62588
rect 9111 62528 9175 62532
rect 9191 62588 9255 62592
rect 9191 62532 9195 62588
rect 9195 62532 9251 62588
rect 9251 62532 9255 62588
rect 9191 62528 9255 62532
rect 9271 62588 9335 62592
rect 9271 62532 9275 62588
rect 9275 62532 9331 62588
rect 9331 62532 9335 62588
rect 9271 62528 9335 62532
rect 9351 62588 9415 62592
rect 9351 62532 9355 62588
rect 9355 62532 9411 62588
rect 9411 62532 9415 62588
rect 9351 62528 9415 62532
rect 4215 62044 4279 62048
rect 4215 61988 4219 62044
rect 4219 61988 4275 62044
rect 4275 61988 4279 62044
rect 4215 61984 4279 61988
rect 4295 62044 4359 62048
rect 4295 61988 4299 62044
rect 4299 61988 4355 62044
rect 4355 61988 4359 62044
rect 4295 61984 4359 61988
rect 4375 62044 4439 62048
rect 4375 61988 4379 62044
rect 4379 61988 4435 62044
rect 4435 61988 4439 62044
rect 4375 61984 4439 61988
rect 4455 62044 4519 62048
rect 4455 61988 4459 62044
rect 4459 61988 4515 62044
rect 4515 61988 4519 62044
rect 4455 61984 4519 61988
rect 7479 62044 7543 62048
rect 7479 61988 7483 62044
rect 7483 61988 7539 62044
rect 7539 61988 7543 62044
rect 7479 61984 7543 61988
rect 7559 62044 7623 62048
rect 7559 61988 7563 62044
rect 7563 61988 7619 62044
rect 7619 61988 7623 62044
rect 7559 61984 7623 61988
rect 7639 62044 7703 62048
rect 7639 61988 7643 62044
rect 7643 61988 7699 62044
rect 7699 61988 7703 62044
rect 7639 61984 7703 61988
rect 7719 62044 7783 62048
rect 7719 61988 7723 62044
rect 7723 61988 7779 62044
rect 7779 61988 7783 62044
rect 7719 61984 7783 61988
rect 2584 61500 2648 61504
rect 2584 61444 2588 61500
rect 2588 61444 2644 61500
rect 2644 61444 2648 61500
rect 2584 61440 2648 61444
rect 2664 61500 2728 61504
rect 2664 61444 2668 61500
rect 2668 61444 2724 61500
rect 2724 61444 2728 61500
rect 2664 61440 2728 61444
rect 2744 61500 2808 61504
rect 2744 61444 2748 61500
rect 2748 61444 2804 61500
rect 2804 61444 2808 61500
rect 2744 61440 2808 61444
rect 2824 61500 2888 61504
rect 2824 61444 2828 61500
rect 2828 61444 2884 61500
rect 2884 61444 2888 61500
rect 2824 61440 2888 61444
rect 5847 61500 5911 61504
rect 5847 61444 5851 61500
rect 5851 61444 5907 61500
rect 5907 61444 5911 61500
rect 5847 61440 5911 61444
rect 5927 61500 5991 61504
rect 5927 61444 5931 61500
rect 5931 61444 5987 61500
rect 5987 61444 5991 61500
rect 5927 61440 5991 61444
rect 6007 61500 6071 61504
rect 6007 61444 6011 61500
rect 6011 61444 6067 61500
rect 6067 61444 6071 61500
rect 6007 61440 6071 61444
rect 6087 61500 6151 61504
rect 6087 61444 6091 61500
rect 6091 61444 6147 61500
rect 6147 61444 6151 61500
rect 6087 61440 6151 61444
rect 9111 61500 9175 61504
rect 9111 61444 9115 61500
rect 9115 61444 9171 61500
rect 9171 61444 9175 61500
rect 9111 61440 9175 61444
rect 9191 61500 9255 61504
rect 9191 61444 9195 61500
rect 9195 61444 9251 61500
rect 9251 61444 9255 61500
rect 9191 61440 9255 61444
rect 9271 61500 9335 61504
rect 9271 61444 9275 61500
rect 9275 61444 9331 61500
rect 9331 61444 9335 61500
rect 9271 61440 9335 61444
rect 9351 61500 9415 61504
rect 9351 61444 9355 61500
rect 9355 61444 9411 61500
rect 9411 61444 9415 61500
rect 9351 61440 9415 61444
rect 4215 60956 4279 60960
rect 4215 60900 4219 60956
rect 4219 60900 4275 60956
rect 4275 60900 4279 60956
rect 4215 60896 4279 60900
rect 4295 60956 4359 60960
rect 4295 60900 4299 60956
rect 4299 60900 4355 60956
rect 4355 60900 4359 60956
rect 4295 60896 4359 60900
rect 4375 60956 4439 60960
rect 4375 60900 4379 60956
rect 4379 60900 4435 60956
rect 4435 60900 4439 60956
rect 4375 60896 4439 60900
rect 4455 60956 4519 60960
rect 4455 60900 4459 60956
rect 4459 60900 4515 60956
rect 4515 60900 4519 60956
rect 4455 60896 4519 60900
rect 7479 60956 7543 60960
rect 7479 60900 7483 60956
rect 7483 60900 7539 60956
rect 7539 60900 7543 60956
rect 7479 60896 7543 60900
rect 7559 60956 7623 60960
rect 7559 60900 7563 60956
rect 7563 60900 7619 60956
rect 7619 60900 7623 60956
rect 7559 60896 7623 60900
rect 7639 60956 7703 60960
rect 7639 60900 7643 60956
rect 7643 60900 7699 60956
rect 7699 60900 7703 60956
rect 7639 60896 7703 60900
rect 7719 60956 7783 60960
rect 7719 60900 7723 60956
rect 7723 60900 7779 60956
rect 7779 60900 7783 60956
rect 7719 60896 7783 60900
rect 2584 60412 2648 60416
rect 2584 60356 2588 60412
rect 2588 60356 2644 60412
rect 2644 60356 2648 60412
rect 2584 60352 2648 60356
rect 2664 60412 2728 60416
rect 2664 60356 2668 60412
rect 2668 60356 2724 60412
rect 2724 60356 2728 60412
rect 2664 60352 2728 60356
rect 2744 60412 2808 60416
rect 2744 60356 2748 60412
rect 2748 60356 2804 60412
rect 2804 60356 2808 60412
rect 2744 60352 2808 60356
rect 2824 60412 2888 60416
rect 2824 60356 2828 60412
rect 2828 60356 2884 60412
rect 2884 60356 2888 60412
rect 2824 60352 2888 60356
rect 5847 60412 5911 60416
rect 5847 60356 5851 60412
rect 5851 60356 5907 60412
rect 5907 60356 5911 60412
rect 5847 60352 5911 60356
rect 5927 60412 5991 60416
rect 5927 60356 5931 60412
rect 5931 60356 5987 60412
rect 5987 60356 5991 60412
rect 5927 60352 5991 60356
rect 6007 60412 6071 60416
rect 6007 60356 6011 60412
rect 6011 60356 6067 60412
rect 6067 60356 6071 60412
rect 6007 60352 6071 60356
rect 6087 60412 6151 60416
rect 6087 60356 6091 60412
rect 6091 60356 6147 60412
rect 6147 60356 6151 60412
rect 6087 60352 6151 60356
rect 9111 60412 9175 60416
rect 9111 60356 9115 60412
rect 9115 60356 9171 60412
rect 9171 60356 9175 60412
rect 9111 60352 9175 60356
rect 9191 60412 9255 60416
rect 9191 60356 9195 60412
rect 9195 60356 9251 60412
rect 9251 60356 9255 60412
rect 9191 60352 9255 60356
rect 9271 60412 9335 60416
rect 9271 60356 9275 60412
rect 9275 60356 9331 60412
rect 9331 60356 9335 60412
rect 9271 60352 9335 60356
rect 9351 60412 9415 60416
rect 9351 60356 9355 60412
rect 9355 60356 9411 60412
rect 9411 60356 9415 60412
rect 9351 60352 9415 60356
rect 4215 59868 4279 59872
rect 4215 59812 4219 59868
rect 4219 59812 4275 59868
rect 4275 59812 4279 59868
rect 4215 59808 4279 59812
rect 4295 59868 4359 59872
rect 4295 59812 4299 59868
rect 4299 59812 4355 59868
rect 4355 59812 4359 59868
rect 4295 59808 4359 59812
rect 4375 59868 4439 59872
rect 4375 59812 4379 59868
rect 4379 59812 4435 59868
rect 4435 59812 4439 59868
rect 4375 59808 4439 59812
rect 4455 59868 4519 59872
rect 4455 59812 4459 59868
rect 4459 59812 4515 59868
rect 4515 59812 4519 59868
rect 4455 59808 4519 59812
rect 7479 59868 7543 59872
rect 7479 59812 7483 59868
rect 7483 59812 7539 59868
rect 7539 59812 7543 59868
rect 7479 59808 7543 59812
rect 7559 59868 7623 59872
rect 7559 59812 7563 59868
rect 7563 59812 7619 59868
rect 7619 59812 7623 59868
rect 7559 59808 7623 59812
rect 7639 59868 7703 59872
rect 7639 59812 7643 59868
rect 7643 59812 7699 59868
rect 7699 59812 7703 59868
rect 7639 59808 7703 59812
rect 7719 59868 7783 59872
rect 7719 59812 7723 59868
rect 7723 59812 7779 59868
rect 7779 59812 7783 59868
rect 7719 59808 7783 59812
rect 2584 59324 2648 59328
rect 2584 59268 2588 59324
rect 2588 59268 2644 59324
rect 2644 59268 2648 59324
rect 2584 59264 2648 59268
rect 2664 59324 2728 59328
rect 2664 59268 2668 59324
rect 2668 59268 2724 59324
rect 2724 59268 2728 59324
rect 2664 59264 2728 59268
rect 2744 59324 2808 59328
rect 2744 59268 2748 59324
rect 2748 59268 2804 59324
rect 2804 59268 2808 59324
rect 2744 59264 2808 59268
rect 2824 59324 2888 59328
rect 2824 59268 2828 59324
rect 2828 59268 2884 59324
rect 2884 59268 2888 59324
rect 2824 59264 2888 59268
rect 5847 59324 5911 59328
rect 5847 59268 5851 59324
rect 5851 59268 5907 59324
rect 5907 59268 5911 59324
rect 5847 59264 5911 59268
rect 5927 59324 5991 59328
rect 5927 59268 5931 59324
rect 5931 59268 5987 59324
rect 5987 59268 5991 59324
rect 5927 59264 5991 59268
rect 6007 59324 6071 59328
rect 6007 59268 6011 59324
rect 6011 59268 6067 59324
rect 6067 59268 6071 59324
rect 6007 59264 6071 59268
rect 6087 59324 6151 59328
rect 6087 59268 6091 59324
rect 6091 59268 6147 59324
rect 6147 59268 6151 59324
rect 6087 59264 6151 59268
rect 9111 59324 9175 59328
rect 9111 59268 9115 59324
rect 9115 59268 9171 59324
rect 9171 59268 9175 59324
rect 9111 59264 9175 59268
rect 9191 59324 9255 59328
rect 9191 59268 9195 59324
rect 9195 59268 9251 59324
rect 9251 59268 9255 59324
rect 9191 59264 9255 59268
rect 9271 59324 9335 59328
rect 9271 59268 9275 59324
rect 9275 59268 9331 59324
rect 9331 59268 9335 59324
rect 9271 59264 9335 59268
rect 9351 59324 9415 59328
rect 9351 59268 9355 59324
rect 9355 59268 9411 59324
rect 9411 59268 9415 59324
rect 9351 59264 9415 59268
rect 4215 58780 4279 58784
rect 4215 58724 4219 58780
rect 4219 58724 4275 58780
rect 4275 58724 4279 58780
rect 4215 58720 4279 58724
rect 4295 58780 4359 58784
rect 4295 58724 4299 58780
rect 4299 58724 4355 58780
rect 4355 58724 4359 58780
rect 4295 58720 4359 58724
rect 4375 58780 4439 58784
rect 4375 58724 4379 58780
rect 4379 58724 4435 58780
rect 4435 58724 4439 58780
rect 4375 58720 4439 58724
rect 4455 58780 4519 58784
rect 4455 58724 4459 58780
rect 4459 58724 4515 58780
rect 4515 58724 4519 58780
rect 4455 58720 4519 58724
rect 7479 58780 7543 58784
rect 7479 58724 7483 58780
rect 7483 58724 7539 58780
rect 7539 58724 7543 58780
rect 7479 58720 7543 58724
rect 7559 58780 7623 58784
rect 7559 58724 7563 58780
rect 7563 58724 7619 58780
rect 7619 58724 7623 58780
rect 7559 58720 7623 58724
rect 7639 58780 7703 58784
rect 7639 58724 7643 58780
rect 7643 58724 7699 58780
rect 7699 58724 7703 58780
rect 7639 58720 7703 58724
rect 7719 58780 7783 58784
rect 7719 58724 7723 58780
rect 7723 58724 7779 58780
rect 7779 58724 7783 58780
rect 7719 58720 7783 58724
rect 2584 58236 2648 58240
rect 2584 58180 2588 58236
rect 2588 58180 2644 58236
rect 2644 58180 2648 58236
rect 2584 58176 2648 58180
rect 2664 58236 2728 58240
rect 2664 58180 2668 58236
rect 2668 58180 2724 58236
rect 2724 58180 2728 58236
rect 2664 58176 2728 58180
rect 2744 58236 2808 58240
rect 2744 58180 2748 58236
rect 2748 58180 2804 58236
rect 2804 58180 2808 58236
rect 2744 58176 2808 58180
rect 2824 58236 2888 58240
rect 2824 58180 2828 58236
rect 2828 58180 2884 58236
rect 2884 58180 2888 58236
rect 2824 58176 2888 58180
rect 5847 58236 5911 58240
rect 5847 58180 5851 58236
rect 5851 58180 5907 58236
rect 5907 58180 5911 58236
rect 5847 58176 5911 58180
rect 5927 58236 5991 58240
rect 5927 58180 5931 58236
rect 5931 58180 5987 58236
rect 5987 58180 5991 58236
rect 5927 58176 5991 58180
rect 6007 58236 6071 58240
rect 6007 58180 6011 58236
rect 6011 58180 6067 58236
rect 6067 58180 6071 58236
rect 6007 58176 6071 58180
rect 6087 58236 6151 58240
rect 6087 58180 6091 58236
rect 6091 58180 6147 58236
rect 6147 58180 6151 58236
rect 6087 58176 6151 58180
rect 9111 58236 9175 58240
rect 9111 58180 9115 58236
rect 9115 58180 9171 58236
rect 9171 58180 9175 58236
rect 9111 58176 9175 58180
rect 9191 58236 9255 58240
rect 9191 58180 9195 58236
rect 9195 58180 9251 58236
rect 9251 58180 9255 58236
rect 9191 58176 9255 58180
rect 9271 58236 9335 58240
rect 9271 58180 9275 58236
rect 9275 58180 9331 58236
rect 9331 58180 9335 58236
rect 9271 58176 9335 58180
rect 9351 58236 9415 58240
rect 9351 58180 9355 58236
rect 9355 58180 9411 58236
rect 9411 58180 9415 58236
rect 9351 58176 9415 58180
rect 4215 57692 4279 57696
rect 4215 57636 4219 57692
rect 4219 57636 4275 57692
rect 4275 57636 4279 57692
rect 4215 57632 4279 57636
rect 4295 57692 4359 57696
rect 4295 57636 4299 57692
rect 4299 57636 4355 57692
rect 4355 57636 4359 57692
rect 4295 57632 4359 57636
rect 4375 57692 4439 57696
rect 4375 57636 4379 57692
rect 4379 57636 4435 57692
rect 4435 57636 4439 57692
rect 4375 57632 4439 57636
rect 4455 57692 4519 57696
rect 4455 57636 4459 57692
rect 4459 57636 4515 57692
rect 4515 57636 4519 57692
rect 4455 57632 4519 57636
rect 7479 57692 7543 57696
rect 7479 57636 7483 57692
rect 7483 57636 7539 57692
rect 7539 57636 7543 57692
rect 7479 57632 7543 57636
rect 7559 57692 7623 57696
rect 7559 57636 7563 57692
rect 7563 57636 7619 57692
rect 7619 57636 7623 57692
rect 7559 57632 7623 57636
rect 7639 57692 7703 57696
rect 7639 57636 7643 57692
rect 7643 57636 7699 57692
rect 7699 57636 7703 57692
rect 7639 57632 7703 57636
rect 7719 57692 7783 57696
rect 7719 57636 7723 57692
rect 7723 57636 7779 57692
rect 7779 57636 7783 57692
rect 7719 57632 7783 57636
rect 3188 57564 3252 57628
rect 2268 57292 2332 57356
rect 2584 57148 2648 57152
rect 2584 57092 2588 57148
rect 2588 57092 2644 57148
rect 2644 57092 2648 57148
rect 2584 57088 2648 57092
rect 2664 57148 2728 57152
rect 2664 57092 2668 57148
rect 2668 57092 2724 57148
rect 2724 57092 2728 57148
rect 2664 57088 2728 57092
rect 2744 57148 2808 57152
rect 2744 57092 2748 57148
rect 2748 57092 2804 57148
rect 2804 57092 2808 57148
rect 2744 57088 2808 57092
rect 2824 57148 2888 57152
rect 2824 57092 2828 57148
rect 2828 57092 2884 57148
rect 2884 57092 2888 57148
rect 2824 57088 2888 57092
rect 5847 57148 5911 57152
rect 5847 57092 5851 57148
rect 5851 57092 5907 57148
rect 5907 57092 5911 57148
rect 5847 57088 5911 57092
rect 5927 57148 5991 57152
rect 5927 57092 5931 57148
rect 5931 57092 5987 57148
rect 5987 57092 5991 57148
rect 5927 57088 5991 57092
rect 6007 57148 6071 57152
rect 6007 57092 6011 57148
rect 6011 57092 6067 57148
rect 6067 57092 6071 57148
rect 6007 57088 6071 57092
rect 6087 57148 6151 57152
rect 6087 57092 6091 57148
rect 6091 57092 6147 57148
rect 6147 57092 6151 57148
rect 6087 57088 6151 57092
rect 9111 57148 9175 57152
rect 9111 57092 9115 57148
rect 9115 57092 9171 57148
rect 9171 57092 9175 57148
rect 9111 57088 9175 57092
rect 9191 57148 9255 57152
rect 9191 57092 9195 57148
rect 9195 57092 9251 57148
rect 9251 57092 9255 57148
rect 9191 57088 9255 57092
rect 9271 57148 9335 57152
rect 9271 57092 9275 57148
rect 9275 57092 9331 57148
rect 9331 57092 9335 57148
rect 9271 57088 9335 57092
rect 9351 57148 9415 57152
rect 9351 57092 9355 57148
rect 9355 57092 9411 57148
rect 9411 57092 9415 57148
rect 9351 57088 9415 57092
rect 4215 56604 4279 56608
rect 4215 56548 4219 56604
rect 4219 56548 4275 56604
rect 4275 56548 4279 56604
rect 4215 56544 4279 56548
rect 4295 56604 4359 56608
rect 4295 56548 4299 56604
rect 4299 56548 4355 56604
rect 4355 56548 4359 56604
rect 4295 56544 4359 56548
rect 4375 56604 4439 56608
rect 4375 56548 4379 56604
rect 4379 56548 4435 56604
rect 4435 56548 4439 56604
rect 4375 56544 4439 56548
rect 4455 56604 4519 56608
rect 4455 56548 4459 56604
rect 4459 56548 4515 56604
rect 4515 56548 4519 56604
rect 4455 56544 4519 56548
rect 7479 56604 7543 56608
rect 7479 56548 7483 56604
rect 7483 56548 7539 56604
rect 7539 56548 7543 56604
rect 7479 56544 7543 56548
rect 7559 56604 7623 56608
rect 7559 56548 7563 56604
rect 7563 56548 7619 56604
rect 7619 56548 7623 56604
rect 7559 56544 7623 56548
rect 7639 56604 7703 56608
rect 7639 56548 7643 56604
rect 7643 56548 7699 56604
rect 7699 56548 7703 56604
rect 7639 56544 7703 56548
rect 7719 56604 7783 56608
rect 7719 56548 7723 56604
rect 7723 56548 7779 56604
rect 7779 56548 7783 56604
rect 7719 56544 7783 56548
rect 3372 56204 3436 56268
rect 2584 56060 2648 56064
rect 2584 56004 2588 56060
rect 2588 56004 2644 56060
rect 2644 56004 2648 56060
rect 2584 56000 2648 56004
rect 2664 56060 2728 56064
rect 2664 56004 2668 56060
rect 2668 56004 2724 56060
rect 2724 56004 2728 56060
rect 2664 56000 2728 56004
rect 2744 56060 2808 56064
rect 2744 56004 2748 56060
rect 2748 56004 2804 56060
rect 2804 56004 2808 56060
rect 2744 56000 2808 56004
rect 2824 56060 2888 56064
rect 2824 56004 2828 56060
rect 2828 56004 2884 56060
rect 2884 56004 2888 56060
rect 2824 56000 2888 56004
rect 5847 56060 5911 56064
rect 5847 56004 5851 56060
rect 5851 56004 5907 56060
rect 5907 56004 5911 56060
rect 5847 56000 5911 56004
rect 5927 56060 5991 56064
rect 5927 56004 5931 56060
rect 5931 56004 5987 56060
rect 5987 56004 5991 56060
rect 5927 56000 5991 56004
rect 6007 56060 6071 56064
rect 6007 56004 6011 56060
rect 6011 56004 6067 56060
rect 6067 56004 6071 56060
rect 6007 56000 6071 56004
rect 6087 56060 6151 56064
rect 6087 56004 6091 56060
rect 6091 56004 6147 56060
rect 6147 56004 6151 56060
rect 6087 56000 6151 56004
rect 9111 56060 9175 56064
rect 9111 56004 9115 56060
rect 9115 56004 9171 56060
rect 9171 56004 9175 56060
rect 9111 56000 9175 56004
rect 9191 56060 9255 56064
rect 9191 56004 9195 56060
rect 9195 56004 9251 56060
rect 9251 56004 9255 56060
rect 9191 56000 9255 56004
rect 9271 56060 9335 56064
rect 9271 56004 9275 56060
rect 9275 56004 9331 56060
rect 9331 56004 9335 56060
rect 9271 56000 9335 56004
rect 9351 56060 9415 56064
rect 9351 56004 9355 56060
rect 9355 56004 9411 56060
rect 9411 56004 9415 56060
rect 9351 56000 9415 56004
rect 4215 55516 4279 55520
rect 4215 55460 4219 55516
rect 4219 55460 4275 55516
rect 4275 55460 4279 55516
rect 4215 55456 4279 55460
rect 4295 55516 4359 55520
rect 4295 55460 4299 55516
rect 4299 55460 4355 55516
rect 4355 55460 4359 55516
rect 4295 55456 4359 55460
rect 4375 55516 4439 55520
rect 4375 55460 4379 55516
rect 4379 55460 4435 55516
rect 4435 55460 4439 55516
rect 4375 55456 4439 55460
rect 4455 55516 4519 55520
rect 4455 55460 4459 55516
rect 4459 55460 4515 55516
rect 4515 55460 4519 55516
rect 4455 55456 4519 55460
rect 7479 55516 7543 55520
rect 7479 55460 7483 55516
rect 7483 55460 7539 55516
rect 7539 55460 7543 55516
rect 7479 55456 7543 55460
rect 7559 55516 7623 55520
rect 7559 55460 7563 55516
rect 7563 55460 7619 55516
rect 7619 55460 7623 55516
rect 7559 55456 7623 55460
rect 7639 55516 7703 55520
rect 7639 55460 7643 55516
rect 7643 55460 7699 55516
rect 7699 55460 7703 55516
rect 7639 55456 7703 55460
rect 7719 55516 7783 55520
rect 7719 55460 7723 55516
rect 7723 55460 7779 55516
rect 7779 55460 7783 55516
rect 7719 55456 7783 55460
rect 3188 55448 3252 55452
rect 3188 55392 3202 55448
rect 3202 55392 3252 55448
rect 3188 55388 3252 55392
rect 2584 54972 2648 54976
rect 2584 54916 2588 54972
rect 2588 54916 2644 54972
rect 2644 54916 2648 54972
rect 2584 54912 2648 54916
rect 2664 54972 2728 54976
rect 2664 54916 2668 54972
rect 2668 54916 2724 54972
rect 2724 54916 2728 54972
rect 2664 54912 2728 54916
rect 2744 54972 2808 54976
rect 2744 54916 2748 54972
rect 2748 54916 2804 54972
rect 2804 54916 2808 54972
rect 2744 54912 2808 54916
rect 2824 54972 2888 54976
rect 2824 54916 2828 54972
rect 2828 54916 2884 54972
rect 2884 54916 2888 54972
rect 2824 54912 2888 54916
rect 5847 54972 5911 54976
rect 5847 54916 5851 54972
rect 5851 54916 5907 54972
rect 5907 54916 5911 54972
rect 5847 54912 5911 54916
rect 5927 54972 5991 54976
rect 5927 54916 5931 54972
rect 5931 54916 5987 54972
rect 5987 54916 5991 54972
rect 5927 54912 5991 54916
rect 6007 54972 6071 54976
rect 6007 54916 6011 54972
rect 6011 54916 6067 54972
rect 6067 54916 6071 54972
rect 6007 54912 6071 54916
rect 6087 54972 6151 54976
rect 6087 54916 6091 54972
rect 6091 54916 6147 54972
rect 6147 54916 6151 54972
rect 6087 54912 6151 54916
rect 9111 54972 9175 54976
rect 9111 54916 9115 54972
rect 9115 54916 9171 54972
rect 9171 54916 9175 54972
rect 9111 54912 9175 54916
rect 9191 54972 9255 54976
rect 9191 54916 9195 54972
rect 9195 54916 9251 54972
rect 9251 54916 9255 54972
rect 9191 54912 9255 54916
rect 9271 54972 9335 54976
rect 9271 54916 9275 54972
rect 9275 54916 9331 54972
rect 9331 54916 9335 54972
rect 9271 54912 9335 54916
rect 9351 54972 9415 54976
rect 9351 54916 9355 54972
rect 9355 54916 9411 54972
rect 9411 54916 9415 54972
rect 9351 54912 9415 54916
rect 1900 54572 1964 54636
rect 4215 54428 4279 54432
rect 4215 54372 4219 54428
rect 4219 54372 4275 54428
rect 4275 54372 4279 54428
rect 4215 54368 4279 54372
rect 4295 54428 4359 54432
rect 4295 54372 4299 54428
rect 4299 54372 4355 54428
rect 4355 54372 4359 54428
rect 4295 54368 4359 54372
rect 4375 54428 4439 54432
rect 4375 54372 4379 54428
rect 4379 54372 4435 54428
rect 4435 54372 4439 54428
rect 4375 54368 4439 54372
rect 4455 54428 4519 54432
rect 4455 54372 4459 54428
rect 4459 54372 4515 54428
rect 4515 54372 4519 54428
rect 4455 54368 4519 54372
rect 7479 54428 7543 54432
rect 7479 54372 7483 54428
rect 7483 54372 7539 54428
rect 7539 54372 7543 54428
rect 7479 54368 7543 54372
rect 7559 54428 7623 54432
rect 7559 54372 7563 54428
rect 7563 54372 7619 54428
rect 7619 54372 7623 54428
rect 7559 54368 7623 54372
rect 7639 54428 7703 54432
rect 7639 54372 7643 54428
rect 7643 54372 7699 54428
rect 7699 54372 7703 54428
rect 7639 54368 7703 54372
rect 7719 54428 7783 54432
rect 7719 54372 7723 54428
rect 7723 54372 7779 54428
rect 7779 54372 7783 54428
rect 7719 54368 7783 54372
rect 2584 53884 2648 53888
rect 2584 53828 2588 53884
rect 2588 53828 2644 53884
rect 2644 53828 2648 53884
rect 2584 53824 2648 53828
rect 2664 53884 2728 53888
rect 2664 53828 2668 53884
rect 2668 53828 2724 53884
rect 2724 53828 2728 53884
rect 2664 53824 2728 53828
rect 2744 53884 2808 53888
rect 2744 53828 2748 53884
rect 2748 53828 2804 53884
rect 2804 53828 2808 53884
rect 2744 53824 2808 53828
rect 2824 53884 2888 53888
rect 2824 53828 2828 53884
rect 2828 53828 2884 53884
rect 2884 53828 2888 53884
rect 2824 53824 2888 53828
rect 5847 53884 5911 53888
rect 5847 53828 5851 53884
rect 5851 53828 5907 53884
rect 5907 53828 5911 53884
rect 5847 53824 5911 53828
rect 5927 53884 5991 53888
rect 5927 53828 5931 53884
rect 5931 53828 5987 53884
rect 5987 53828 5991 53884
rect 5927 53824 5991 53828
rect 6007 53884 6071 53888
rect 6007 53828 6011 53884
rect 6011 53828 6067 53884
rect 6067 53828 6071 53884
rect 6007 53824 6071 53828
rect 6087 53884 6151 53888
rect 6087 53828 6091 53884
rect 6091 53828 6147 53884
rect 6147 53828 6151 53884
rect 6087 53824 6151 53828
rect 9111 53884 9175 53888
rect 9111 53828 9115 53884
rect 9115 53828 9171 53884
rect 9171 53828 9175 53884
rect 9111 53824 9175 53828
rect 9191 53884 9255 53888
rect 9191 53828 9195 53884
rect 9195 53828 9251 53884
rect 9251 53828 9255 53884
rect 9191 53824 9255 53828
rect 9271 53884 9335 53888
rect 9271 53828 9275 53884
rect 9275 53828 9331 53884
rect 9331 53828 9335 53884
rect 9271 53824 9335 53828
rect 9351 53884 9415 53888
rect 9351 53828 9355 53884
rect 9355 53828 9411 53884
rect 9411 53828 9415 53884
rect 9351 53824 9415 53828
rect 4215 53340 4279 53344
rect 4215 53284 4219 53340
rect 4219 53284 4275 53340
rect 4275 53284 4279 53340
rect 4215 53280 4279 53284
rect 4295 53340 4359 53344
rect 4295 53284 4299 53340
rect 4299 53284 4355 53340
rect 4355 53284 4359 53340
rect 4295 53280 4359 53284
rect 4375 53340 4439 53344
rect 4375 53284 4379 53340
rect 4379 53284 4435 53340
rect 4435 53284 4439 53340
rect 4375 53280 4439 53284
rect 4455 53340 4519 53344
rect 4455 53284 4459 53340
rect 4459 53284 4515 53340
rect 4515 53284 4519 53340
rect 4455 53280 4519 53284
rect 7479 53340 7543 53344
rect 7479 53284 7483 53340
rect 7483 53284 7539 53340
rect 7539 53284 7543 53340
rect 7479 53280 7543 53284
rect 7559 53340 7623 53344
rect 7559 53284 7563 53340
rect 7563 53284 7619 53340
rect 7619 53284 7623 53340
rect 7559 53280 7623 53284
rect 7639 53340 7703 53344
rect 7639 53284 7643 53340
rect 7643 53284 7699 53340
rect 7699 53284 7703 53340
rect 7639 53280 7703 53284
rect 7719 53340 7783 53344
rect 7719 53284 7723 53340
rect 7723 53284 7779 53340
rect 7779 53284 7783 53340
rect 7719 53280 7783 53284
rect 2584 52796 2648 52800
rect 2584 52740 2588 52796
rect 2588 52740 2644 52796
rect 2644 52740 2648 52796
rect 2584 52736 2648 52740
rect 2664 52796 2728 52800
rect 2664 52740 2668 52796
rect 2668 52740 2724 52796
rect 2724 52740 2728 52796
rect 2664 52736 2728 52740
rect 2744 52796 2808 52800
rect 2744 52740 2748 52796
rect 2748 52740 2804 52796
rect 2804 52740 2808 52796
rect 2744 52736 2808 52740
rect 2824 52796 2888 52800
rect 2824 52740 2828 52796
rect 2828 52740 2884 52796
rect 2884 52740 2888 52796
rect 2824 52736 2888 52740
rect 5847 52796 5911 52800
rect 5847 52740 5851 52796
rect 5851 52740 5907 52796
rect 5907 52740 5911 52796
rect 5847 52736 5911 52740
rect 5927 52796 5991 52800
rect 5927 52740 5931 52796
rect 5931 52740 5987 52796
rect 5987 52740 5991 52796
rect 5927 52736 5991 52740
rect 6007 52796 6071 52800
rect 6007 52740 6011 52796
rect 6011 52740 6067 52796
rect 6067 52740 6071 52796
rect 6007 52736 6071 52740
rect 6087 52796 6151 52800
rect 6087 52740 6091 52796
rect 6091 52740 6147 52796
rect 6147 52740 6151 52796
rect 6087 52736 6151 52740
rect 9111 52796 9175 52800
rect 9111 52740 9115 52796
rect 9115 52740 9171 52796
rect 9171 52740 9175 52796
rect 9111 52736 9175 52740
rect 9191 52796 9255 52800
rect 9191 52740 9195 52796
rect 9195 52740 9251 52796
rect 9251 52740 9255 52796
rect 9191 52736 9255 52740
rect 9271 52796 9335 52800
rect 9271 52740 9275 52796
rect 9275 52740 9331 52796
rect 9331 52740 9335 52796
rect 9271 52736 9335 52740
rect 9351 52796 9415 52800
rect 9351 52740 9355 52796
rect 9355 52740 9411 52796
rect 9411 52740 9415 52796
rect 9351 52736 9415 52740
rect 4215 52252 4279 52256
rect 4215 52196 4219 52252
rect 4219 52196 4275 52252
rect 4275 52196 4279 52252
rect 4215 52192 4279 52196
rect 4295 52252 4359 52256
rect 4295 52196 4299 52252
rect 4299 52196 4355 52252
rect 4355 52196 4359 52252
rect 4295 52192 4359 52196
rect 4375 52252 4439 52256
rect 4375 52196 4379 52252
rect 4379 52196 4435 52252
rect 4435 52196 4439 52252
rect 4375 52192 4439 52196
rect 4455 52252 4519 52256
rect 4455 52196 4459 52252
rect 4459 52196 4515 52252
rect 4515 52196 4519 52252
rect 4455 52192 4519 52196
rect 7479 52252 7543 52256
rect 7479 52196 7483 52252
rect 7483 52196 7539 52252
rect 7539 52196 7543 52252
rect 7479 52192 7543 52196
rect 7559 52252 7623 52256
rect 7559 52196 7563 52252
rect 7563 52196 7619 52252
rect 7619 52196 7623 52252
rect 7559 52192 7623 52196
rect 7639 52252 7703 52256
rect 7639 52196 7643 52252
rect 7643 52196 7699 52252
rect 7699 52196 7703 52252
rect 7639 52192 7703 52196
rect 7719 52252 7783 52256
rect 7719 52196 7723 52252
rect 7723 52196 7779 52252
rect 7779 52196 7783 52252
rect 7719 52192 7783 52196
rect 2584 51708 2648 51712
rect 2584 51652 2588 51708
rect 2588 51652 2644 51708
rect 2644 51652 2648 51708
rect 2584 51648 2648 51652
rect 2664 51708 2728 51712
rect 2664 51652 2668 51708
rect 2668 51652 2724 51708
rect 2724 51652 2728 51708
rect 2664 51648 2728 51652
rect 2744 51708 2808 51712
rect 2744 51652 2748 51708
rect 2748 51652 2804 51708
rect 2804 51652 2808 51708
rect 2744 51648 2808 51652
rect 2824 51708 2888 51712
rect 2824 51652 2828 51708
rect 2828 51652 2884 51708
rect 2884 51652 2888 51708
rect 2824 51648 2888 51652
rect 5847 51708 5911 51712
rect 5847 51652 5851 51708
rect 5851 51652 5907 51708
rect 5907 51652 5911 51708
rect 5847 51648 5911 51652
rect 5927 51708 5991 51712
rect 5927 51652 5931 51708
rect 5931 51652 5987 51708
rect 5987 51652 5991 51708
rect 5927 51648 5991 51652
rect 6007 51708 6071 51712
rect 6007 51652 6011 51708
rect 6011 51652 6067 51708
rect 6067 51652 6071 51708
rect 6007 51648 6071 51652
rect 6087 51708 6151 51712
rect 6087 51652 6091 51708
rect 6091 51652 6147 51708
rect 6147 51652 6151 51708
rect 6087 51648 6151 51652
rect 9111 51708 9175 51712
rect 9111 51652 9115 51708
rect 9115 51652 9171 51708
rect 9171 51652 9175 51708
rect 9111 51648 9175 51652
rect 9191 51708 9255 51712
rect 9191 51652 9195 51708
rect 9195 51652 9251 51708
rect 9251 51652 9255 51708
rect 9191 51648 9255 51652
rect 9271 51708 9335 51712
rect 9271 51652 9275 51708
rect 9275 51652 9331 51708
rect 9331 51652 9335 51708
rect 9271 51648 9335 51652
rect 9351 51708 9415 51712
rect 9351 51652 9355 51708
rect 9355 51652 9411 51708
rect 9411 51652 9415 51708
rect 9351 51648 9415 51652
rect 3924 51172 3988 51236
rect 4215 51164 4279 51168
rect 4215 51108 4219 51164
rect 4219 51108 4275 51164
rect 4275 51108 4279 51164
rect 4215 51104 4279 51108
rect 4295 51164 4359 51168
rect 4295 51108 4299 51164
rect 4299 51108 4355 51164
rect 4355 51108 4359 51164
rect 4295 51104 4359 51108
rect 4375 51164 4439 51168
rect 4375 51108 4379 51164
rect 4379 51108 4435 51164
rect 4435 51108 4439 51164
rect 4375 51104 4439 51108
rect 4455 51164 4519 51168
rect 4455 51108 4459 51164
rect 4459 51108 4515 51164
rect 4515 51108 4519 51164
rect 4455 51104 4519 51108
rect 7479 51164 7543 51168
rect 7479 51108 7483 51164
rect 7483 51108 7539 51164
rect 7539 51108 7543 51164
rect 7479 51104 7543 51108
rect 7559 51164 7623 51168
rect 7559 51108 7563 51164
rect 7563 51108 7619 51164
rect 7619 51108 7623 51164
rect 7559 51104 7623 51108
rect 7639 51164 7703 51168
rect 7639 51108 7643 51164
rect 7643 51108 7699 51164
rect 7699 51108 7703 51164
rect 7639 51104 7703 51108
rect 7719 51164 7783 51168
rect 7719 51108 7723 51164
rect 7723 51108 7779 51164
rect 7779 51108 7783 51164
rect 7719 51104 7783 51108
rect 2084 51036 2148 51100
rect 3740 51096 3804 51100
rect 3740 51040 3754 51096
rect 3754 51040 3804 51096
rect 3740 51036 3804 51040
rect 6316 50900 6380 50964
rect 2268 50764 2332 50828
rect 3004 50764 3068 50828
rect 3372 50824 3436 50828
rect 3372 50768 3386 50824
rect 3386 50768 3436 50824
rect 3372 50764 3436 50768
rect 1900 50628 1964 50692
rect 2584 50620 2648 50624
rect 2584 50564 2588 50620
rect 2588 50564 2644 50620
rect 2644 50564 2648 50620
rect 2584 50560 2648 50564
rect 2664 50620 2728 50624
rect 2664 50564 2668 50620
rect 2668 50564 2724 50620
rect 2724 50564 2728 50620
rect 2664 50560 2728 50564
rect 2744 50620 2808 50624
rect 2744 50564 2748 50620
rect 2748 50564 2804 50620
rect 2804 50564 2808 50620
rect 2744 50560 2808 50564
rect 2824 50620 2888 50624
rect 2824 50564 2828 50620
rect 2828 50564 2884 50620
rect 2884 50564 2888 50620
rect 2824 50560 2888 50564
rect 5847 50620 5911 50624
rect 5847 50564 5851 50620
rect 5851 50564 5907 50620
rect 5907 50564 5911 50620
rect 5847 50560 5911 50564
rect 5927 50620 5991 50624
rect 5927 50564 5931 50620
rect 5931 50564 5987 50620
rect 5987 50564 5991 50620
rect 5927 50560 5991 50564
rect 6007 50620 6071 50624
rect 6007 50564 6011 50620
rect 6011 50564 6067 50620
rect 6067 50564 6071 50620
rect 6007 50560 6071 50564
rect 6087 50620 6151 50624
rect 6087 50564 6091 50620
rect 6091 50564 6147 50620
rect 6147 50564 6151 50620
rect 6087 50560 6151 50564
rect 9111 50620 9175 50624
rect 9111 50564 9115 50620
rect 9115 50564 9171 50620
rect 9171 50564 9175 50620
rect 9111 50560 9175 50564
rect 9191 50620 9255 50624
rect 9191 50564 9195 50620
rect 9195 50564 9251 50620
rect 9251 50564 9255 50620
rect 9191 50560 9255 50564
rect 9271 50620 9335 50624
rect 9271 50564 9275 50620
rect 9275 50564 9331 50620
rect 9331 50564 9335 50620
rect 9271 50560 9335 50564
rect 9351 50620 9415 50624
rect 9351 50564 9355 50620
rect 9355 50564 9411 50620
rect 9411 50564 9415 50620
rect 9351 50560 9415 50564
rect 3188 50492 3252 50556
rect 4215 50076 4279 50080
rect 4215 50020 4219 50076
rect 4219 50020 4275 50076
rect 4275 50020 4279 50076
rect 4215 50016 4279 50020
rect 4295 50076 4359 50080
rect 4295 50020 4299 50076
rect 4299 50020 4355 50076
rect 4355 50020 4359 50076
rect 4295 50016 4359 50020
rect 4375 50076 4439 50080
rect 4375 50020 4379 50076
rect 4379 50020 4435 50076
rect 4435 50020 4439 50076
rect 4375 50016 4439 50020
rect 4455 50076 4519 50080
rect 4455 50020 4459 50076
rect 4459 50020 4515 50076
rect 4515 50020 4519 50076
rect 4455 50016 4519 50020
rect 7479 50076 7543 50080
rect 7479 50020 7483 50076
rect 7483 50020 7539 50076
rect 7539 50020 7543 50076
rect 7479 50016 7543 50020
rect 7559 50076 7623 50080
rect 7559 50020 7563 50076
rect 7563 50020 7619 50076
rect 7619 50020 7623 50076
rect 7559 50016 7623 50020
rect 7639 50076 7703 50080
rect 7639 50020 7643 50076
rect 7643 50020 7699 50076
rect 7699 50020 7703 50076
rect 7639 50016 7703 50020
rect 7719 50076 7783 50080
rect 7719 50020 7723 50076
rect 7723 50020 7779 50076
rect 7779 50020 7783 50076
rect 7719 50016 7783 50020
rect 3924 49812 3988 49876
rect 6500 49676 6564 49740
rect 3740 49540 3804 49604
rect 4660 49540 4724 49604
rect 2584 49532 2648 49536
rect 2584 49476 2588 49532
rect 2588 49476 2644 49532
rect 2644 49476 2648 49532
rect 2584 49472 2648 49476
rect 2664 49532 2728 49536
rect 2664 49476 2668 49532
rect 2668 49476 2724 49532
rect 2724 49476 2728 49532
rect 2664 49472 2728 49476
rect 2744 49532 2808 49536
rect 2744 49476 2748 49532
rect 2748 49476 2804 49532
rect 2804 49476 2808 49532
rect 2744 49472 2808 49476
rect 2824 49532 2888 49536
rect 2824 49476 2828 49532
rect 2828 49476 2884 49532
rect 2884 49476 2888 49532
rect 2824 49472 2888 49476
rect 5847 49532 5911 49536
rect 5847 49476 5851 49532
rect 5851 49476 5907 49532
rect 5907 49476 5911 49532
rect 5847 49472 5911 49476
rect 5927 49532 5991 49536
rect 5927 49476 5931 49532
rect 5931 49476 5987 49532
rect 5987 49476 5991 49532
rect 5927 49472 5991 49476
rect 6007 49532 6071 49536
rect 6007 49476 6011 49532
rect 6011 49476 6067 49532
rect 6067 49476 6071 49532
rect 6007 49472 6071 49476
rect 6087 49532 6151 49536
rect 6087 49476 6091 49532
rect 6091 49476 6147 49532
rect 6147 49476 6151 49532
rect 6087 49472 6151 49476
rect 9111 49532 9175 49536
rect 9111 49476 9115 49532
rect 9115 49476 9171 49532
rect 9171 49476 9175 49532
rect 9111 49472 9175 49476
rect 9191 49532 9255 49536
rect 9191 49476 9195 49532
rect 9195 49476 9251 49532
rect 9251 49476 9255 49532
rect 9191 49472 9255 49476
rect 9271 49532 9335 49536
rect 9271 49476 9275 49532
rect 9275 49476 9331 49532
rect 9331 49476 9335 49532
rect 9271 49472 9335 49476
rect 9351 49532 9415 49536
rect 9351 49476 9355 49532
rect 9355 49476 9411 49532
rect 9411 49476 9415 49532
rect 9351 49472 9415 49476
rect 2084 48996 2148 49060
rect 5396 48996 5460 49060
rect 4215 48988 4279 48992
rect 4215 48932 4219 48988
rect 4219 48932 4275 48988
rect 4275 48932 4279 48988
rect 4215 48928 4279 48932
rect 4295 48988 4359 48992
rect 4295 48932 4299 48988
rect 4299 48932 4355 48988
rect 4355 48932 4359 48988
rect 4295 48928 4359 48932
rect 4375 48988 4439 48992
rect 4375 48932 4379 48988
rect 4379 48932 4435 48988
rect 4435 48932 4439 48988
rect 4375 48928 4439 48932
rect 4455 48988 4519 48992
rect 4455 48932 4459 48988
rect 4459 48932 4515 48988
rect 4515 48932 4519 48988
rect 4455 48928 4519 48932
rect 7479 48988 7543 48992
rect 7479 48932 7483 48988
rect 7483 48932 7539 48988
rect 7539 48932 7543 48988
rect 7479 48928 7543 48932
rect 7559 48988 7623 48992
rect 7559 48932 7563 48988
rect 7563 48932 7619 48988
rect 7619 48932 7623 48988
rect 7559 48928 7623 48932
rect 7639 48988 7703 48992
rect 7639 48932 7643 48988
rect 7643 48932 7699 48988
rect 7699 48932 7703 48988
rect 7639 48928 7703 48932
rect 7719 48988 7783 48992
rect 7719 48932 7723 48988
rect 7723 48932 7779 48988
rect 7779 48932 7783 48988
rect 7719 48928 7783 48932
rect 5580 48920 5644 48924
rect 5580 48864 5594 48920
rect 5594 48864 5644 48920
rect 5580 48860 5644 48864
rect 5396 48452 5460 48516
rect 2584 48444 2648 48448
rect 2584 48388 2588 48444
rect 2588 48388 2644 48444
rect 2644 48388 2648 48444
rect 2584 48384 2648 48388
rect 2664 48444 2728 48448
rect 2664 48388 2668 48444
rect 2668 48388 2724 48444
rect 2724 48388 2728 48444
rect 2664 48384 2728 48388
rect 2744 48444 2808 48448
rect 2744 48388 2748 48444
rect 2748 48388 2804 48444
rect 2804 48388 2808 48444
rect 2744 48384 2808 48388
rect 2824 48444 2888 48448
rect 2824 48388 2828 48444
rect 2828 48388 2884 48444
rect 2884 48388 2888 48444
rect 2824 48384 2888 48388
rect 5847 48444 5911 48448
rect 5847 48388 5851 48444
rect 5851 48388 5907 48444
rect 5907 48388 5911 48444
rect 5847 48384 5911 48388
rect 5927 48444 5991 48448
rect 5927 48388 5931 48444
rect 5931 48388 5987 48444
rect 5987 48388 5991 48444
rect 5927 48384 5991 48388
rect 6007 48444 6071 48448
rect 6007 48388 6011 48444
rect 6011 48388 6067 48444
rect 6067 48388 6071 48444
rect 6007 48384 6071 48388
rect 6087 48444 6151 48448
rect 6087 48388 6091 48444
rect 6091 48388 6147 48444
rect 6147 48388 6151 48444
rect 6087 48384 6151 48388
rect 9111 48444 9175 48448
rect 9111 48388 9115 48444
rect 9115 48388 9171 48444
rect 9171 48388 9175 48444
rect 9111 48384 9175 48388
rect 9191 48444 9255 48448
rect 9191 48388 9195 48444
rect 9195 48388 9251 48444
rect 9251 48388 9255 48444
rect 9191 48384 9255 48388
rect 9271 48444 9335 48448
rect 9271 48388 9275 48444
rect 9275 48388 9331 48444
rect 9331 48388 9335 48444
rect 9271 48384 9335 48388
rect 9351 48444 9415 48448
rect 9351 48388 9355 48444
rect 9355 48388 9411 48444
rect 9411 48388 9415 48444
rect 9351 48384 9415 48388
rect 5580 48342 5644 48380
rect 5580 48316 5594 48342
rect 5594 48316 5644 48342
rect 2268 48180 2332 48244
rect 4215 47900 4279 47904
rect 4215 47844 4219 47900
rect 4219 47844 4275 47900
rect 4275 47844 4279 47900
rect 4215 47840 4279 47844
rect 4295 47900 4359 47904
rect 4295 47844 4299 47900
rect 4299 47844 4355 47900
rect 4355 47844 4359 47900
rect 4295 47840 4359 47844
rect 4375 47900 4439 47904
rect 4375 47844 4379 47900
rect 4379 47844 4435 47900
rect 4435 47844 4439 47900
rect 4375 47840 4439 47844
rect 4455 47900 4519 47904
rect 4455 47844 4459 47900
rect 4459 47844 4515 47900
rect 4515 47844 4519 47900
rect 4455 47840 4519 47844
rect 7479 47900 7543 47904
rect 7479 47844 7483 47900
rect 7483 47844 7539 47900
rect 7539 47844 7543 47900
rect 7479 47840 7543 47844
rect 7559 47900 7623 47904
rect 7559 47844 7563 47900
rect 7563 47844 7619 47900
rect 7619 47844 7623 47900
rect 7559 47840 7623 47844
rect 7639 47900 7703 47904
rect 7639 47844 7643 47900
rect 7643 47844 7699 47900
rect 7699 47844 7703 47900
rect 7639 47840 7703 47844
rect 7719 47900 7783 47904
rect 7719 47844 7723 47900
rect 7723 47844 7779 47900
rect 7779 47844 7783 47900
rect 7719 47840 7783 47844
rect 4844 47772 4908 47836
rect 2584 47356 2648 47360
rect 2584 47300 2588 47356
rect 2588 47300 2644 47356
rect 2644 47300 2648 47356
rect 2584 47296 2648 47300
rect 2664 47356 2728 47360
rect 2664 47300 2668 47356
rect 2668 47300 2724 47356
rect 2724 47300 2728 47356
rect 2664 47296 2728 47300
rect 2744 47356 2808 47360
rect 2744 47300 2748 47356
rect 2748 47300 2804 47356
rect 2804 47300 2808 47356
rect 2744 47296 2808 47300
rect 2824 47356 2888 47360
rect 2824 47300 2828 47356
rect 2828 47300 2884 47356
rect 2884 47300 2888 47356
rect 2824 47296 2888 47300
rect 5847 47356 5911 47360
rect 5847 47300 5851 47356
rect 5851 47300 5907 47356
rect 5907 47300 5911 47356
rect 5847 47296 5911 47300
rect 5927 47356 5991 47360
rect 5927 47300 5931 47356
rect 5931 47300 5987 47356
rect 5987 47300 5991 47356
rect 5927 47296 5991 47300
rect 6007 47356 6071 47360
rect 6007 47300 6011 47356
rect 6011 47300 6067 47356
rect 6067 47300 6071 47356
rect 6007 47296 6071 47300
rect 6087 47356 6151 47360
rect 6087 47300 6091 47356
rect 6091 47300 6147 47356
rect 6147 47300 6151 47356
rect 6087 47296 6151 47300
rect 9111 47356 9175 47360
rect 9111 47300 9115 47356
rect 9115 47300 9171 47356
rect 9171 47300 9175 47356
rect 9111 47296 9175 47300
rect 9191 47356 9255 47360
rect 9191 47300 9195 47356
rect 9195 47300 9251 47356
rect 9251 47300 9255 47356
rect 9191 47296 9255 47300
rect 9271 47356 9335 47360
rect 9271 47300 9275 47356
rect 9275 47300 9331 47356
rect 9331 47300 9335 47356
rect 9271 47296 9335 47300
rect 9351 47356 9415 47360
rect 9351 47300 9355 47356
rect 9355 47300 9411 47356
rect 9411 47300 9415 47356
rect 9351 47296 9415 47300
rect 4215 46812 4279 46816
rect 4215 46756 4219 46812
rect 4219 46756 4275 46812
rect 4275 46756 4279 46812
rect 4215 46752 4279 46756
rect 4295 46812 4359 46816
rect 4295 46756 4299 46812
rect 4299 46756 4355 46812
rect 4355 46756 4359 46812
rect 4295 46752 4359 46756
rect 4375 46812 4439 46816
rect 4375 46756 4379 46812
rect 4379 46756 4435 46812
rect 4435 46756 4439 46812
rect 4375 46752 4439 46756
rect 4455 46812 4519 46816
rect 4455 46756 4459 46812
rect 4459 46756 4515 46812
rect 4515 46756 4519 46812
rect 4455 46752 4519 46756
rect 7479 46812 7543 46816
rect 7479 46756 7483 46812
rect 7483 46756 7539 46812
rect 7539 46756 7543 46812
rect 7479 46752 7543 46756
rect 7559 46812 7623 46816
rect 7559 46756 7563 46812
rect 7563 46756 7619 46812
rect 7619 46756 7623 46812
rect 7559 46752 7623 46756
rect 7639 46812 7703 46816
rect 7639 46756 7643 46812
rect 7643 46756 7699 46812
rect 7699 46756 7703 46812
rect 7639 46752 7703 46756
rect 7719 46812 7783 46816
rect 7719 46756 7723 46812
rect 7723 46756 7779 46812
rect 7779 46756 7783 46812
rect 7719 46752 7783 46756
rect 3188 46684 3252 46748
rect 3924 46412 3988 46476
rect 2584 46268 2648 46272
rect 2584 46212 2588 46268
rect 2588 46212 2644 46268
rect 2644 46212 2648 46268
rect 2584 46208 2648 46212
rect 2664 46268 2728 46272
rect 2664 46212 2668 46268
rect 2668 46212 2724 46268
rect 2724 46212 2728 46268
rect 2664 46208 2728 46212
rect 2744 46268 2808 46272
rect 2744 46212 2748 46268
rect 2748 46212 2804 46268
rect 2804 46212 2808 46268
rect 2744 46208 2808 46212
rect 2824 46268 2888 46272
rect 2824 46212 2828 46268
rect 2828 46212 2884 46268
rect 2884 46212 2888 46268
rect 2824 46208 2888 46212
rect 5847 46268 5911 46272
rect 5847 46212 5851 46268
rect 5851 46212 5907 46268
rect 5907 46212 5911 46268
rect 5847 46208 5911 46212
rect 5927 46268 5991 46272
rect 5927 46212 5931 46268
rect 5931 46212 5987 46268
rect 5987 46212 5991 46268
rect 5927 46208 5991 46212
rect 6007 46268 6071 46272
rect 6007 46212 6011 46268
rect 6011 46212 6067 46268
rect 6067 46212 6071 46268
rect 6007 46208 6071 46212
rect 6087 46268 6151 46272
rect 6087 46212 6091 46268
rect 6091 46212 6147 46268
rect 6147 46212 6151 46268
rect 6087 46208 6151 46212
rect 5028 46140 5092 46204
rect 3004 46004 3068 46068
rect 9111 46268 9175 46272
rect 9111 46212 9115 46268
rect 9115 46212 9171 46268
rect 9171 46212 9175 46268
rect 9111 46208 9175 46212
rect 9191 46268 9255 46272
rect 9191 46212 9195 46268
rect 9195 46212 9251 46268
rect 9251 46212 9255 46268
rect 9191 46208 9255 46212
rect 9271 46268 9335 46272
rect 9271 46212 9275 46268
rect 9275 46212 9331 46268
rect 9331 46212 9335 46268
rect 9271 46208 9335 46212
rect 9351 46268 9415 46272
rect 9351 46212 9355 46268
rect 9355 46212 9411 46268
rect 9411 46212 9415 46268
rect 9351 46208 9415 46212
rect 4215 45724 4279 45728
rect 4215 45668 4219 45724
rect 4219 45668 4275 45724
rect 4275 45668 4279 45724
rect 4215 45664 4279 45668
rect 4295 45724 4359 45728
rect 4295 45668 4299 45724
rect 4299 45668 4355 45724
rect 4355 45668 4359 45724
rect 4295 45664 4359 45668
rect 4375 45724 4439 45728
rect 4375 45668 4379 45724
rect 4379 45668 4435 45724
rect 4435 45668 4439 45724
rect 4375 45664 4439 45668
rect 4455 45724 4519 45728
rect 4455 45668 4459 45724
rect 4459 45668 4515 45724
rect 4515 45668 4519 45724
rect 4455 45664 4519 45668
rect 7479 45724 7543 45728
rect 7479 45668 7483 45724
rect 7483 45668 7539 45724
rect 7539 45668 7543 45724
rect 7479 45664 7543 45668
rect 7559 45724 7623 45728
rect 7559 45668 7563 45724
rect 7563 45668 7619 45724
rect 7619 45668 7623 45724
rect 7559 45664 7623 45668
rect 7639 45724 7703 45728
rect 7639 45668 7643 45724
rect 7643 45668 7699 45724
rect 7699 45668 7703 45724
rect 7639 45664 7703 45668
rect 7719 45724 7783 45728
rect 7719 45668 7723 45724
rect 7723 45668 7779 45724
rect 7779 45668 7783 45724
rect 7719 45664 7783 45668
rect 2584 45180 2648 45184
rect 2584 45124 2588 45180
rect 2588 45124 2644 45180
rect 2644 45124 2648 45180
rect 2584 45120 2648 45124
rect 2664 45180 2728 45184
rect 2664 45124 2668 45180
rect 2668 45124 2724 45180
rect 2724 45124 2728 45180
rect 2664 45120 2728 45124
rect 2744 45180 2808 45184
rect 2744 45124 2748 45180
rect 2748 45124 2804 45180
rect 2804 45124 2808 45180
rect 2744 45120 2808 45124
rect 2824 45180 2888 45184
rect 2824 45124 2828 45180
rect 2828 45124 2884 45180
rect 2884 45124 2888 45180
rect 2824 45120 2888 45124
rect 5847 45180 5911 45184
rect 5847 45124 5851 45180
rect 5851 45124 5907 45180
rect 5907 45124 5911 45180
rect 5847 45120 5911 45124
rect 5927 45180 5991 45184
rect 5927 45124 5931 45180
rect 5931 45124 5987 45180
rect 5987 45124 5991 45180
rect 5927 45120 5991 45124
rect 6007 45180 6071 45184
rect 6007 45124 6011 45180
rect 6011 45124 6067 45180
rect 6067 45124 6071 45180
rect 6007 45120 6071 45124
rect 6087 45180 6151 45184
rect 6087 45124 6091 45180
rect 6091 45124 6147 45180
rect 6147 45124 6151 45180
rect 6087 45120 6151 45124
rect 9111 45180 9175 45184
rect 9111 45124 9115 45180
rect 9115 45124 9171 45180
rect 9171 45124 9175 45180
rect 9111 45120 9175 45124
rect 9191 45180 9255 45184
rect 9191 45124 9195 45180
rect 9195 45124 9251 45180
rect 9251 45124 9255 45180
rect 9191 45120 9255 45124
rect 9271 45180 9335 45184
rect 9271 45124 9275 45180
rect 9275 45124 9331 45180
rect 9331 45124 9335 45180
rect 9271 45120 9335 45124
rect 9351 45180 9415 45184
rect 9351 45124 9355 45180
rect 9355 45124 9411 45180
rect 9411 45124 9415 45180
rect 9351 45120 9415 45124
rect 2084 45112 2148 45116
rect 2084 45056 2098 45112
rect 2098 45056 2148 45112
rect 2084 45052 2148 45056
rect 3004 45052 3068 45116
rect 4215 44636 4279 44640
rect 4215 44580 4219 44636
rect 4219 44580 4275 44636
rect 4275 44580 4279 44636
rect 4215 44576 4279 44580
rect 4295 44636 4359 44640
rect 4295 44580 4299 44636
rect 4299 44580 4355 44636
rect 4355 44580 4359 44636
rect 4295 44576 4359 44580
rect 4375 44636 4439 44640
rect 4375 44580 4379 44636
rect 4379 44580 4435 44636
rect 4435 44580 4439 44636
rect 4375 44576 4439 44580
rect 4455 44636 4519 44640
rect 4455 44580 4459 44636
rect 4459 44580 4515 44636
rect 4515 44580 4519 44636
rect 4455 44576 4519 44580
rect 7479 44636 7543 44640
rect 7479 44580 7483 44636
rect 7483 44580 7539 44636
rect 7539 44580 7543 44636
rect 7479 44576 7543 44580
rect 7559 44636 7623 44640
rect 7559 44580 7563 44636
rect 7563 44580 7619 44636
rect 7619 44580 7623 44636
rect 7559 44576 7623 44580
rect 7639 44636 7703 44640
rect 7639 44580 7643 44636
rect 7643 44580 7699 44636
rect 7699 44580 7703 44636
rect 7639 44576 7703 44580
rect 7719 44636 7783 44640
rect 7719 44580 7723 44636
rect 7723 44580 7779 44636
rect 7779 44580 7783 44636
rect 7719 44576 7783 44580
rect 2584 44092 2648 44096
rect 2584 44036 2588 44092
rect 2588 44036 2644 44092
rect 2644 44036 2648 44092
rect 2584 44032 2648 44036
rect 2664 44092 2728 44096
rect 2664 44036 2668 44092
rect 2668 44036 2724 44092
rect 2724 44036 2728 44092
rect 2664 44032 2728 44036
rect 2744 44092 2808 44096
rect 2744 44036 2748 44092
rect 2748 44036 2804 44092
rect 2804 44036 2808 44092
rect 2744 44032 2808 44036
rect 2824 44092 2888 44096
rect 2824 44036 2828 44092
rect 2828 44036 2884 44092
rect 2884 44036 2888 44092
rect 2824 44032 2888 44036
rect 5847 44092 5911 44096
rect 5847 44036 5851 44092
rect 5851 44036 5907 44092
rect 5907 44036 5911 44092
rect 5847 44032 5911 44036
rect 5927 44092 5991 44096
rect 5927 44036 5931 44092
rect 5931 44036 5987 44092
rect 5987 44036 5991 44092
rect 5927 44032 5991 44036
rect 6007 44092 6071 44096
rect 6007 44036 6011 44092
rect 6011 44036 6067 44092
rect 6067 44036 6071 44092
rect 6007 44032 6071 44036
rect 6087 44092 6151 44096
rect 6087 44036 6091 44092
rect 6091 44036 6147 44092
rect 6147 44036 6151 44092
rect 6087 44032 6151 44036
rect 9111 44092 9175 44096
rect 9111 44036 9115 44092
rect 9115 44036 9171 44092
rect 9171 44036 9175 44092
rect 9111 44032 9175 44036
rect 9191 44092 9255 44096
rect 9191 44036 9195 44092
rect 9195 44036 9251 44092
rect 9251 44036 9255 44092
rect 9191 44032 9255 44036
rect 9271 44092 9335 44096
rect 9271 44036 9275 44092
rect 9275 44036 9331 44092
rect 9331 44036 9335 44092
rect 9271 44032 9335 44036
rect 9351 44092 9415 44096
rect 9351 44036 9355 44092
rect 9355 44036 9411 44092
rect 9411 44036 9415 44092
rect 9351 44032 9415 44036
rect 4215 43548 4279 43552
rect 4215 43492 4219 43548
rect 4219 43492 4275 43548
rect 4275 43492 4279 43548
rect 4215 43488 4279 43492
rect 4295 43548 4359 43552
rect 4295 43492 4299 43548
rect 4299 43492 4355 43548
rect 4355 43492 4359 43548
rect 4295 43488 4359 43492
rect 4375 43548 4439 43552
rect 4375 43492 4379 43548
rect 4379 43492 4435 43548
rect 4435 43492 4439 43548
rect 4375 43488 4439 43492
rect 4455 43548 4519 43552
rect 4455 43492 4459 43548
rect 4459 43492 4515 43548
rect 4515 43492 4519 43548
rect 4455 43488 4519 43492
rect 7479 43548 7543 43552
rect 7479 43492 7483 43548
rect 7483 43492 7539 43548
rect 7539 43492 7543 43548
rect 7479 43488 7543 43492
rect 7559 43548 7623 43552
rect 7559 43492 7563 43548
rect 7563 43492 7619 43548
rect 7619 43492 7623 43548
rect 7559 43488 7623 43492
rect 7639 43548 7703 43552
rect 7639 43492 7643 43548
rect 7643 43492 7699 43548
rect 7699 43492 7703 43548
rect 7639 43488 7703 43492
rect 7719 43548 7783 43552
rect 7719 43492 7723 43548
rect 7723 43492 7779 43548
rect 7779 43492 7783 43548
rect 7719 43488 7783 43492
rect 2268 43480 2332 43484
rect 2268 43424 2318 43480
rect 2318 43424 2332 43480
rect 2268 43420 2332 43424
rect 3188 43284 3252 43348
rect 4660 43284 4724 43348
rect 2584 43004 2648 43008
rect 2584 42948 2588 43004
rect 2588 42948 2644 43004
rect 2644 42948 2648 43004
rect 2584 42944 2648 42948
rect 2664 43004 2728 43008
rect 2664 42948 2668 43004
rect 2668 42948 2724 43004
rect 2724 42948 2728 43004
rect 2664 42944 2728 42948
rect 2744 43004 2808 43008
rect 2744 42948 2748 43004
rect 2748 42948 2804 43004
rect 2804 42948 2808 43004
rect 2744 42944 2808 42948
rect 2824 43004 2888 43008
rect 2824 42948 2828 43004
rect 2828 42948 2884 43004
rect 2884 42948 2888 43004
rect 2824 42944 2888 42948
rect 5847 43004 5911 43008
rect 5847 42948 5851 43004
rect 5851 42948 5907 43004
rect 5907 42948 5911 43004
rect 5847 42944 5911 42948
rect 5927 43004 5991 43008
rect 5927 42948 5931 43004
rect 5931 42948 5987 43004
rect 5987 42948 5991 43004
rect 5927 42944 5991 42948
rect 6007 43004 6071 43008
rect 6007 42948 6011 43004
rect 6011 42948 6067 43004
rect 6067 42948 6071 43004
rect 6007 42944 6071 42948
rect 6087 43004 6151 43008
rect 6087 42948 6091 43004
rect 6091 42948 6147 43004
rect 6147 42948 6151 43004
rect 6087 42944 6151 42948
rect 9111 43004 9175 43008
rect 9111 42948 9115 43004
rect 9115 42948 9171 43004
rect 9171 42948 9175 43004
rect 9111 42944 9175 42948
rect 9191 43004 9255 43008
rect 9191 42948 9195 43004
rect 9195 42948 9251 43004
rect 9251 42948 9255 43004
rect 9191 42944 9255 42948
rect 9271 43004 9335 43008
rect 9271 42948 9275 43004
rect 9275 42948 9331 43004
rect 9331 42948 9335 43004
rect 9271 42944 9335 42948
rect 9351 43004 9415 43008
rect 9351 42948 9355 43004
rect 9355 42948 9411 43004
rect 9411 42948 9415 43004
rect 9351 42944 9415 42948
rect 4215 42460 4279 42464
rect 4215 42404 4219 42460
rect 4219 42404 4275 42460
rect 4275 42404 4279 42460
rect 4215 42400 4279 42404
rect 4295 42460 4359 42464
rect 4295 42404 4299 42460
rect 4299 42404 4355 42460
rect 4355 42404 4359 42460
rect 4295 42400 4359 42404
rect 4375 42460 4439 42464
rect 4375 42404 4379 42460
rect 4379 42404 4435 42460
rect 4435 42404 4439 42460
rect 4375 42400 4439 42404
rect 4455 42460 4519 42464
rect 4455 42404 4459 42460
rect 4459 42404 4515 42460
rect 4515 42404 4519 42460
rect 4455 42400 4519 42404
rect 7479 42460 7543 42464
rect 7479 42404 7483 42460
rect 7483 42404 7539 42460
rect 7539 42404 7543 42460
rect 7479 42400 7543 42404
rect 7559 42460 7623 42464
rect 7559 42404 7563 42460
rect 7563 42404 7619 42460
rect 7619 42404 7623 42460
rect 7559 42400 7623 42404
rect 7639 42460 7703 42464
rect 7639 42404 7643 42460
rect 7643 42404 7699 42460
rect 7699 42404 7703 42460
rect 7639 42400 7703 42404
rect 7719 42460 7783 42464
rect 7719 42404 7723 42460
rect 7723 42404 7779 42460
rect 7779 42404 7783 42460
rect 7719 42400 7783 42404
rect 4844 42196 4908 42260
rect 2084 42120 2148 42124
rect 2084 42064 2098 42120
rect 2098 42064 2148 42120
rect 2084 42060 2148 42064
rect 5028 41984 5092 41988
rect 5028 41928 5078 41984
rect 5078 41928 5092 41984
rect 5028 41924 5092 41928
rect 2584 41916 2648 41920
rect 2584 41860 2588 41916
rect 2588 41860 2644 41916
rect 2644 41860 2648 41916
rect 2584 41856 2648 41860
rect 2664 41916 2728 41920
rect 2664 41860 2668 41916
rect 2668 41860 2724 41916
rect 2724 41860 2728 41916
rect 2664 41856 2728 41860
rect 2744 41916 2808 41920
rect 2744 41860 2748 41916
rect 2748 41860 2804 41916
rect 2804 41860 2808 41916
rect 2744 41856 2808 41860
rect 2824 41916 2888 41920
rect 2824 41860 2828 41916
rect 2828 41860 2884 41916
rect 2884 41860 2888 41916
rect 2824 41856 2888 41860
rect 5847 41916 5911 41920
rect 5847 41860 5851 41916
rect 5851 41860 5907 41916
rect 5907 41860 5911 41916
rect 5847 41856 5911 41860
rect 5927 41916 5991 41920
rect 5927 41860 5931 41916
rect 5931 41860 5987 41916
rect 5987 41860 5991 41916
rect 5927 41856 5991 41860
rect 6007 41916 6071 41920
rect 6007 41860 6011 41916
rect 6011 41860 6067 41916
rect 6067 41860 6071 41916
rect 6007 41856 6071 41860
rect 6087 41916 6151 41920
rect 6087 41860 6091 41916
rect 6091 41860 6147 41916
rect 6147 41860 6151 41916
rect 6087 41856 6151 41860
rect 9111 41916 9175 41920
rect 9111 41860 9115 41916
rect 9115 41860 9171 41916
rect 9171 41860 9175 41916
rect 9111 41856 9175 41860
rect 9191 41916 9255 41920
rect 9191 41860 9195 41916
rect 9195 41860 9251 41916
rect 9251 41860 9255 41916
rect 9191 41856 9255 41860
rect 9271 41916 9335 41920
rect 9271 41860 9275 41916
rect 9275 41860 9331 41916
rect 9331 41860 9335 41916
rect 9271 41856 9335 41860
rect 9351 41916 9415 41920
rect 9351 41860 9355 41916
rect 9355 41860 9411 41916
rect 9411 41860 9415 41916
rect 9351 41856 9415 41860
rect 5396 41652 5460 41716
rect 5212 41516 5276 41580
rect 6316 41516 6380 41580
rect 4215 41372 4279 41376
rect 4215 41316 4219 41372
rect 4219 41316 4275 41372
rect 4275 41316 4279 41372
rect 4215 41312 4279 41316
rect 4295 41372 4359 41376
rect 4295 41316 4299 41372
rect 4299 41316 4355 41372
rect 4355 41316 4359 41372
rect 4295 41312 4359 41316
rect 4375 41372 4439 41376
rect 4375 41316 4379 41372
rect 4379 41316 4435 41372
rect 4435 41316 4439 41372
rect 4375 41312 4439 41316
rect 4455 41372 4519 41376
rect 4455 41316 4459 41372
rect 4459 41316 4515 41372
rect 4515 41316 4519 41372
rect 4455 41312 4519 41316
rect 7479 41372 7543 41376
rect 7479 41316 7483 41372
rect 7483 41316 7539 41372
rect 7539 41316 7543 41372
rect 7479 41312 7543 41316
rect 7559 41372 7623 41376
rect 7559 41316 7563 41372
rect 7563 41316 7619 41372
rect 7619 41316 7623 41372
rect 7559 41312 7623 41316
rect 7639 41372 7703 41376
rect 7639 41316 7643 41372
rect 7643 41316 7699 41372
rect 7699 41316 7703 41372
rect 7639 41312 7703 41316
rect 7719 41372 7783 41376
rect 7719 41316 7723 41372
rect 7723 41316 7779 41372
rect 7779 41316 7783 41372
rect 7719 41312 7783 41316
rect 2268 41304 2332 41308
rect 2268 41248 2318 41304
rect 2318 41248 2332 41304
rect 2268 41244 2332 41248
rect 6500 41244 6564 41308
rect 1164 41108 1228 41172
rect 2584 40828 2648 40832
rect 2584 40772 2588 40828
rect 2588 40772 2644 40828
rect 2644 40772 2648 40828
rect 2584 40768 2648 40772
rect 2664 40828 2728 40832
rect 2664 40772 2668 40828
rect 2668 40772 2724 40828
rect 2724 40772 2728 40828
rect 2664 40768 2728 40772
rect 2744 40828 2808 40832
rect 2744 40772 2748 40828
rect 2748 40772 2804 40828
rect 2804 40772 2808 40828
rect 2744 40768 2808 40772
rect 2824 40828 2888 40832
rect 2824 40772 2828 40828
rect 2828 40772 2884 40828
rect 2884 40772 2888 40828
rect 2824 40768 2888 40772
rect 5847 40828 5911 40832
rect 5847 40772 5851 40828
rect 5851 40772 5907 40828
rect 5907 40772 5911 40828
rect 5847 40768 5911 40772
rect 5927 40828 5991 40832
rect 5927 40772 5931 40828
rect 5931 40772 5987 40828
rect 5987 40772 5991 40828
rect 5927 40768 5991 40772
rect 6007 40828 6071 40832
rect 6007 40772 6011 40828
rect 6011 40772 6067 40828
rect 6067 40772 6071 40828
rect 6007 40768 6071 40772
rect 6087 40828 6151 40832
rect 6087 40772 6091 40828
rect 6091 40772 6147 40828
rect 6147 40772 6151 40828
rect 6087 40768 6151 40772
rect 9111 40828 9175 40832
rect 9111 40772 9115 40828
rect 9115 40772 9171 40828
rect 9171 40772 9175 40828
rect 9111 40768 9175 40772
rect 9191 40828 9255 40832
rect 9191 40772 9195 40828
rect 9195 40772 9251 40828
rect 9251 40772 9255 40828
rect 9191 40768 9255 40772
rect 9271 40828 9335 40832
rect 9271 40772 9275 40828
rect 9275 40772 9331 40828
rect 9331 40772 9335 40828
rect 9271 40768 9335 40772
rect 9351 40828 9415 40832
rect 9351 40772 9355 40828
rect 9355 40772 9411 40828
rect 9411 40772 9415 40828
rect 9351 40768 9415 40772
rect 4215 40284 4279 40288
rect 4215 40228 4219 40284
rect 4219 40228 4275 40284
rect 4275 40228 4279 40284
rect 4215 40224 4279 40228
rect 4295 40284 4359 40288
rect 4295 40228 4299 40284
rect 4299 40228 4355 40284
rect 4355 40228 4359 40284
rect 4295 40224 4359 40228
rect 4375 40284 4439 40288
rect 4375 40228 4379 40284
rect 4379 40228 4435 40284
rect 4435 40228 4439 40284
rect 4375 40224 4439 40228
rect 4455 40284 4519 40288
rect 4455 40228 4459 40284
rect 4459 40228 4515 40284
rect 4515 40228 4519 40284
rect 4455 40224 4519 40228
rect 7479 40284 7543 40288
rect 7479 40228 7483 40284
rect 7483 40228 7539 40284
rect 7539 40228 7543 40284
rect 7479 40224 7543 40228
rect 7559 40284 7623 40288
rect 7559 40228 7563 40284
rect 7563 40228 7619 40284
rect 7619 40228 7623 40284
rect 7559 40224 7623 40228
rect 7639 40284 7703 40288
rect 7639 40228 7643 40284
rect 7643 40228 7699 40284
rect 7699 40228 7703 40284
rect 7639 40224 7703 40228
rect 7719 40284 7783 40288
rect 7719 40228 7723 40284
rect 7723 40228 7779 40284
rect 7779 40228 7783 40284
rect 7719 40224 7783 40228
rect 5212 39808 5276 39812
rect 5212 39752 5226 39808
rect 5226 39752 5276 39808
rect 5212 39748 5276 39752
rect 2584 39740 2648 39744
rect 2584 39684 2588 39740
rect 2588 39684 2644 39740
rect 2644 39684 2648 39740
rect 2584 39680 2648 39684
rect 2664 39740 2728 39744
rect 2664 39684 2668 39740
rect 2668 39684 2724 39740
rect 2724 39684 2728 39740
rect 2664 39680 2728 39684
rect 2744 39740 2808 39744
rect 2744 39684 2748 39740
rect 2748 39684 2804 39740
rect 2804 39684 2808 39740
rect 2744 39680 2808 39684
rect 2824 39740 2888 39744
rect 2824 39684 2828 39740
rect 2828 39684 2884 39740
rect 2884 39684 2888 39740
rect 2824 39680 2888 39684
rect 5847 39740 5911 39744
rect 5847 39684 5851 39740
rect 5851 39684 5907 39740
rect 5907 39684 5911 39740
rect 5847 39680 5911 39684
rect 5927 39740 5991 39744
rect 5927 39684 5931 39740
rect 5931 39684 5987 39740
rect 5987 39684 5991 39740
rect 5927 39680 5991 39684
rect 6007 39740 6071 39744
rect 6007 39684 6011 39740
rect 6011 39684 6067 39740
rect 6067 39684 6071 39740
rect 6007 39680 6071 39684
rect 6087 39740 6151 39744
rect 6087 39684 6091 39740
rect 6091 39684 6147 39740
rect 6147 39684 6151 39740
rect 6087 39680 6151 39684
rect 9111 39740 9175 39744
rect 9111 39684 9115 39740
rect 9115 39684 9171 39740
rect 9171 39684 9175 39740
rect 9111 39680 9175 39684
rect 9191 39740 9255 39744
rect 9191 39684 9195 39740
rect 9195 39684 9251 39740
rect 9251 39684 9255 39740
rect 9191 39680 9255 39684
rect 9271 39740 9335 39744
rect 9271 39684 9275 39740
rect 9275 39684 9331 39740
rect 9331 39684 9335 39740
rect 9271 39680 9335 39684
rect 9351 39740 9415 39744
rect 9351 39684 9355 39740
rect 9355 39684 9411 39740
rect 9411 39684 9415 39740
rect 9351 39680 9415 39684
rect 5396 39476 5460 39540
rect 4215 39196 4279 39200
rect 4215 39140 4219 39196
rect 4219 39140 4275 39196
rect 4275 39140 4279 39196
rect 4215 39136 4279 39140
rect 4295 39196 4359 39200
rect 4295 39140 4299 39196
rect 4299 39140 4355 39196
rect 4355 39140 4359 39196
rect 4295 39136 4359 39140
rect 4375 39196 4439 39200
rect 4375 39140 4379 39196
rect 4379 39140 4435 39196
rect 4435 39140 4439 39196
rect 4375 39136 4439 39140
rect 4455 39196 4519 39200
rect 4455 39140 4459 39196
rect 4459 39140 4515 39196
rect 4515 39140 4519 39196
rect 4455 39136 4519 39140
rect 7479 39196 7543 39200
rect 7479 39140 7483 39196
rect 7483 39140 7539 39196
rect 7539 39140 7543 39196
rect 7479 39136 7543 39140
rect 7559 39196 7623 39200
rect 7559 39140 7563 39196
rect 7563 39140 7619 39196
rect 7619 39140 7623 39196
rect 7559 39136 7623 39140
rect 7639 39196 7703 39200
rect 7639 39140 7643 39196
rect 7643 39140 7699 39196
rect 7699 39140 7703 39196
rect 7639 39136 7703 39140
rect 7719 39196 7783 39200
rect 7719 39140 7723 39196
rect 7723 39140 7779 39196
rect 7779 39140 7783 39196
rect 7719 39136 7783 39140
rect 3924 38796 3988 38860
rect 2084 38660 2148 38724
rect 3004 38720 3068 38724
rect 3004 38664 3018 38720
rect 3018 38664 3068 38720
rect 3004 38660 3068 38664
rect 2584 38652 2648 38656
rect 2584 38596 2588 38652
rect 2588 38596 2644 38652
rect 2644 38596 2648 38652
rect 2584 38592 2648 38596
rect 2664 38652 2728 38656
rect 2664 38596 2668 38652
rect 2668 38596 2724 38652
rect 2724 38596 2728 38652
rect 2664 38592 2728 38596
rect 2744 38652 2808 38656
rect 2744 38596 2748 38652
rect 2748 38596 2804 38652
rect 2804 38596 2808 38652
rect 2744 38592 2808 38596
rect 2824 38652 2888 38656
rect 2824 38596 2828 38652
rect 2828 38596 2884 38652
rect 2884 38596 2888 38652
rect 2824 38592 2888 38596
rect 5847 38652 5911 38656
rect 5847 38596 5851 38652
rect 5851 38596 5907 38652
rect 5907 38596 5911 38652
rect 5847 38592 5911 38596
rect 5927 38652 5991 38656
rect 5927 38596 5931 38652
rect 5931 38596 5987 38652
rect 5987 38596 5991 38652
rect 5927 38592 5991 38596
rect 6007 38652 6071 38656
rect 6007 38596 6011 38652
rect 6011 38596 6067 38652
rect 6067 38596 6071 38652
rect 6007 38592 6071 38596
rect 6087 38652 6151 38656
rect 6087 38596 6091 38652
rect 6091 38596 6147 38652
rect 6147 38596 6151 38652
rect 6087 38592 6151 38596
rect 9111 38652 9175 38656
rect 9111 38596 9115 38652
rect 9115 38596 9171 38652
rect 9171 38596 9175 38652
rect 9111 38592 9175 38596
rect 9191 38652 9255 38656
rect 9191 38596 9195 38652
rect 9195 38596 9251 38652
rect 9251 38596 9255 38652
rect 9191 38592 9255 38596
rect 9271 38652 9335 38656
rect 9271 38596 9275 38652
rect 9275 38596 9331 38652
rect 9331 38596 9335 38652
rect 9271 38592 9335 38596
rect 9351 38652 9415 38656
rect 9351 38596 9355 38652
rect 9355 38596 9411 38652
rect 9411 38596 9415 38652
rect 9351 38592 9415 38596
rect 4215 38108 4279 38112
rect 4215 38052 4219 38108
rect 4219 38052 4275 38108
rect 4275 38052 4279 38108
rect 4215 38048 4279 38052
rect 4295 38108 4359 38112
rect 4295 38052 4299 38108
rect 4299 38052 4355 38108
rect 4355 38052 4359 38108
rect 4295 38048 4359 38052
rect 4375 38108 4439 38112
rect 4375 38052 4379 38108
rect 4379 38052 4435 38108
rect 4435 38052 4439 38108
rect 4375 38048 4439 38052
rect 4455 38108 4519 38112
rect 4455 38052 4459 38108
rect 4459 38052 4515 38108
rect 4515 38052 4519 38108
rect 4455 38048 4519 38052
rect 7479 38108 7543 38112
rect 7479 38052 7483 38108
rect 7483 38052 7539 38108
rect 7539 38052 7543 38108
rect 7479 38048 7543 38052
rect 7559 38108 7623 38112
rect 7559 38052 7563 38108
rect 7563 38052 7619 38108
rect 7619 38052 7623 38108
rect 7559 38048 7623 38052
rect 7639 38108 7703 38112
rect 7639 38052 7643 38108
rect 7643 38052 7699 38108
rect 7699 38052 7703 38108
rect 7639 38048 7703 38052
rect 7719 38108 7783 38112
rect 7719 38052 7723 38108
rect 7723 38052 7779 38108
rect 7779 38052 7783 38108
rect 7719 38048 7783 38052
rect 2584 37564 2648 37568
rect 2584 37508 2588 37564
rect 2588 37508 2644 37564
rect 2644 37508 2648 37564
rect 2584 37504 2648 37508
rect 2664 37564 2728 37568
rect 2664 37508 2668 37564
rect 2668 37508 2724 37564
rect 2724 37508 2728 37564
rect 2664 37504 2728 37508
rect 2744 37564 2808 37568
rect 2744 37508 2748 37564
rect 2748 37508 2804 37564
rect 2804 37508 2808 37564
rect 2744 37504 2808 37508
rect 2824 37564 2888 37568
rect 2824 37508 2828 37564
rect 2828 37508 2884 37564
rect 2884 37508 2888 37564
rect 2824 37504 2888 37508
rect 5847 37564 5911 37568
rect 5847 37508 5851 37564
rect 5851 37508 5907 37564
rect 5907 37508 5911 37564
rect 5847 37504 5911 37508
rect 5927 37564 5991 37568
rect 5927 37508 5931 37564
rect 5931 37508 5987 37564
rect 5987 37508 5991 37564
rect 5927 37504 5991 37508
rect 6007 37564 6071 37568
rect 6007 37508 6011 37564
rect 6011 37508 6067 37564
rect 6067 37508 6071 37564
rect 6007 37504 6071 37508
rect 6087 37564 6151 37568
rect 6087 37508 6091 37564
rect 6091 37508 6147 37564
rect 6147 37508 6151 37564
rect 6087 37504 6151 37508
rect 9111 37564 9175 37568
rect 9111 37508 9115 37564
rect 9115 37508 9171 37564
rect 9171 37508 9175 37564
rect 9111 37504 9175 37508
rect 9191 37564 9255 37568
rect 9191 37508 9195 37564
rect 9195 37508 9251 37564
rect 9251 37508 9255 37564
rect 9191 37504 9255 37508
rect 9271 37564 9335 37568
rect 9271 37508 9275 37564
rect 9275 37508 9331 37564
rect 9331 37508 9335 37564
rect 9271 37504 9335 37508
rect 9351 37564 9415 37568
rect 9351 37508 9355 37564
rect 9355 37508 9411 37564
rect 9411 37508 9415 37564
rect 9351 37504 9415 37508
rect 3740 37300 3804 37364
rect 3004 37224 3068 37228
rect 3004 37168 3018 37224
rect 3018 37168 3068 37224
rect 3004 37164 3068 37168
rect 4215 37020 4279 37024
rect 4215 36964 4219 37020
rect 4219 36964 4275 37020
rect 4275 36964 4279 37020
rect 4215 36960 4279 36964
rect 4295 37020 4359 37024
rect 4295 36964 4299 37020
rect 4299 36964 4355 37020
rect 4355 36964 4359 37020
rect 4295 36960 4359 36964
rect 4375 37020 4439 37024
rect 4375 36964 4379 37020
rect 4379 36964 4435 37020
rect 4435 36964 4439 37020
rect 4375 36960 4439 36964
rect 4455 37020 4519 37024
rect 4455 36964 4459 37020
rect 4459 36964 4515 37020
rect 4515 36964 4519 37020
rect 4455 36960 4519 36964
rect 7479 37020 7543 37024
rect 7479 36964 7483 37020
rect 7483 36964 7539 37020
rect 7539 36964 7543 37020
rect 7479 36960 7543 36964
rect 7559 37020 7623 37024
rect 7559 36964 7563 37020
rect 7563 36964 7619 37020
rect 7619 36964 7623 37020
rect 7559 36960 7623 36964
rect 7639 37020 7703 37024
rect 7639 36964 7643 37020
rect 7643 36964 7699 37020
rect 7699 36964 7703 37020
rect 7639 36960 7703 36964
rect 7719 37020 7783 37024
rect 7719 36964 7723 37020
rect 7723 36964 7779 37020
rect 7779 36964 7783 37020
rect 7719 36960 7783 36964
rect 3556 36680 3620 36684
rect 3556 36624 3570 36680
rect 3570 36624 3620 36680
rect 3556 36620 3620 36624
rect 2584 36476 2648 36480
rect 2584 36420 2588 36476
rect 2588 36420 2644 36476
rect 2644 36420 2648 36476
rect 2584 36416 2648 36420
rect 2664 36476 2728 36480
rect 2664 36420 2668 36476
rect 2668 36420 2724 36476
rect 2724 36420 2728 36476
rect 2664 36416 2728 36420
rect 2744 36476 2808 36480
rect 2744 36420 2748 36476
rect 2748 36420 2804 36476
rect 2804 36420 2808 36476
rect 2744 36416 2808 36420
rect 2824 36476 2888 36480
rect 2824 36420 2828 36476
rect 2828 36420 2884 36476
rect 2884 36420 2888 36476
rect 2824 36416 2888 36420
rect 5847 36476 5911 36480
rect 5847 36420 5851 36476
rect 5851 36420 5907 36476
rect 5907 36420 5911 36476
rect 5847 36416 5911 36420
rect 5927 36476 5991 36480
rect 5927 36420 5931 36476
rect 5931 36420 5987 36476
rect 5987 36420 5991 36476
rect 5927 36416 5991 36420
rect 6007 36476 6071 36480
rect 6007 36420 6011 36476
rect 6011 36420 6067 36476
rect 6067 36420 6071 36476
rect 6007 36416 6071 36420
rect 6087 36476 6151 36480
rect 6087 36420 6091 36476
rect 6091 36420 6147 36476
rect 6147 36420 6151 36476
rect 6087 36416 6151 36420
rect 9111 36476 9175 36480
rect 9111 36420 9115 36476
rect 9115 36420 9171 36476
rect 9171 36420 9175 36476
rect 9111 36416 9175 36420
rect 9191 36476 9255 36480
rect 9191 36420 9195 36476
rect 9195 36420 9251 36476
rect 9251 36420 9255 36476
rect 9191 36416 9255 36420
rect 9271 36476 9335 36480
rect 9271 36420 9275 36476
rect 9275 36420 9331 36476
rect 9331 36420 9335 36476
rect 9271 36416 9335 36420
rect 9351 36476 9415 36480
rect 9351 36420 9355 36476
rect 9355 36420 9411 36476
rect 9411 36420 9415 36476
rect 9351 36416 9415 36420
rect 1532 36136 1596 36140
rect 1532 36080 1546 36136
rect 1546 36080 1596 36136
rect 1532 36076 1596 36080
rect 4215 35932 4279 35936
rect 4215 35876 4219 35932
rect 4219 35876 4275 35932
rect 4275 35876 4279 35932
rect 4215 35872 4279 35876
rect 4295 35932 4359 35936
rect 4295 35876 4299 35932
rect 4299 35876 4355 35932
rect 4355 35876 4359 35932
rect 4295 35872 4359 35876
rect 4375 35932 4439 35936
rect 4375 35876 4379 35932
rect 4379 35876 4435 35932
rect 4435 35876 4439 35932
rect 4375 35872 4439 35876
rect 4455 35932 4519 35936
rect 4455 35876 4459 35932
rect 4459 35876 4515 35932
rect 4515 35876 4519 35932
rect 4455 35872 4519 35876
rect 7479 35932 7543 35936
rect 7479 35876 7483 35932
rect 7483 35876 7539 35932
rect 7539 35876 7543 35932
rect 7479 35872 7543 35876
rect 7559 35932 7623 35936
rect 7559 35876 7563 35932
rect 7563 35876 7619 35932
rect 7619 35876 7623 35932
rect 7559 35872 7623 35876
rect 7639 35932 7703 35936
rect 7639 35876 7643 35932
rect 7643 35876 7699 35932
rect 7699 35876 7703 35932
rect 7639 35872 7703 35876
rect 7719 35932 7783 35936
rect 7719 35876 7723 35932
rect 7723 35876 7779 35932
rect 7779 35876 7783 35932
rect 7719 35872 7783 35876
rect 3740 35456 3804 35460
rect 3740 35400 3754 35456
rect 3754 35400 3804 35456
rect 3740 35396 3804 35400
rect 2584 35388 2648 35392
rect 2584 35332 2588 35388
rect 2588 35332 2644 35388
rect 2644 35332 2648 35388
rect 2584 35328 2648 35332
rect 2664 35388 2728 35392
rect 2664 35332 2668 35388
rect 2668 35332 2724 35388
rect 2724 35332 2728 35388
rect 2664 35328 2728 35332
rect 2744 35388 2808 35392
rect 2744 35332 2748 35388
rect 2748 35332 2804 35388
rect 2804 35332 2808 35388
rect 2744 35328 2808 35332
rect 2824 35388 2888 35392
rect 2824 35332 2828 35388
rect 2828 35332 2884 35388
rect 2884 35332 2888 35388
rect 2824 35328 2888 35332
rect 5847 35388 5911 35392
rect 5847 35332 5851 35388
rect 5851 35332 5907 35388
rect 5907 35332 5911 35388
rect 5847 35328 5911 35332
rect 5927 35388 5991 35392
rect 5927 35332 5931 35388
rect 5931 35332 5987 35388
rect 5987 35332 5991 35388
rect 5927 35328 5991 35332
rect 6007 35388 6071 35392
rect 6007 35332 6011 35388
rect 6011 35332 6067 35388
rect 6067 35332 6071 35388
rect 6007 35328 6071 35332
rect 6087 35388 6151 35392
rect 6087 35332 6091 35388
rect 6091 35332 6147 35388
rect 6147 35332 6151 35388
rect 6087 35328 6151 35332
rect 9111 35388 9175 35392
rect 9111 35332 9115 35388
rect 9115 35332 9171 35388
rect 9171 35332 9175 35388
rect 9111 35328 9175 35332
rect 9191 35388 9255 35392
rect 9191 35332 9195 35388
rect 9195 35332 9251 35388
rect 9251 35332 9255 35388
rect 9191 35328 9255 35332
rect 9271 35388 9335 35392
rect 9271 35332 9275 35388
rect 9275 35332 9331 35388
rect 9331 35332 9335 35388
rect 9271 35328 9335 35332
rect 9351 35388 9415 35392
rect 9351 35332 9355 35388
rect 9355 35332 9411 35388
rect 9411 35332 9415 35388
rect 9351 35328 9415 35332
rect 4215 34844 4279 34848
rect 4215 34788 4219 34844
rect 4219 34788 4275 34844
rect 4275 34788 4279 34844
rect 4215 34784 4279 34788
rect 4295 34844 4359 34848
rect 4295 34788 4299 34844
rect 4299 34788 4355 34844
rect 4355 34788 4359 34844
rect 4295 34784 4359 34788
rect 4375 34844 4439 34848
rect 4375 34788 4379 34844
rect 4379 34788 4435 34844
rect 4435 34788 4439 34844
rect 4375 34784 4439 34788
rect 4455 34844 4519 34848
rect 4455 34788 4459 34844
rect 4459 34788 4515 34844
rect 4515 34788 4519 34844
rect 4455 34784 4519 34788
rect 7479 34844 7543 34848
rect 7479 34788 7483 34844
rect 7483 34788 7539 34844
rect 7539 34788 7543 34844
rect 7479 34784 7543 34788
rect 7559 34844 7623 34848
rect 7559 34788 7563 34844
rect 7563 34788 7619 34844
rect 7619 34788 7623 34844
rect 7559 34784 7623 34788
rect 7639 34844 7703 34848
rect 7639 34788 7643 34844
rect 7643 34788 7699 34844
rect 7699 34788 7703 34844
rect 7639 34784 7703 34788
rect 7719 34844 7783 34848
rect 7719 34788 7723 34844
rect 7723 34788 7779 34844
rect 7779 34788 7783 34844
rect 7719 34784 7783 34788
rect 2584 34300 2648 34304
rect 2584 34244 2588 34300
rect 2588 34244 2644 34300
rect 2644 34244 2648 34300
rect 2584 34240 2648 34244
rect 2664 34300 2728 34304
rect 2664 34244 2668 34300
rect 2668 34244 2724 34300
rect 2724 34244 2728 34300
rect 2664 34240 2728 34244
rect 2744 34300 2808 34304
rect 2744 34244 2748 34300
rect 2748 34244 2804 34300
rect 2804 34244 2808 34300
rect 2744 34240 2808 34244
rect 2824 34300 2888 34304
rect 2824 34244 2828 34300
rect 2828 34244 2884 34300
rect 2884 34244 2888 34300
rect 2824 34240 2888 34244
rect 5847 34300 5911 34304
rect 5847 34244 5851 34300
rect 5851 34244 5907 34300
rect 5907 34244 5911 34300
rect 5847 34240 5911 34244
rect 5927 34300 5991 34304
rect 5927 34244 5931 34300
rect 5931 34244 5987 34300
rect 5987 34244 5991 34300
rect 5927 34240 5991 34244
rect 6007 34300 6071 34304
rect 6007 34244 6011 34300
rect 6011 34244 6067 34300
rect 6067 34244 6071 34300
rect 6007 34240 6071 34244
rect 6087 34300 6151 34304
rect 6087 34244 6091 34300
rect 6091 34244 6147 34300
rect 6147 34244 6151 34300
rect 6087 34240 6151 34244
rect 9111 34300 9175 34304
rect 9111 34244 9115 34300
rect 9115 34244 9171 34300
rect 9171 34244 9175 34300
rect 9111 34240 9175 34244
rect 9191 34300 9255 34304
rect 9191 34244 9195 34300
rect 9195 34244 9251 34300
rect 9251 34244 9255 34300
rect 9191 34240 9255 34244
rect 9271 34300 9335 34304
rect 9271 34244 9275 34300
rect 9275 34244 9331 34300
rect 9331 34244 9335 34300
rect 9271 34240 9335 34244
rect 9351 34300 9415 34304
rect 9351 34244 9355 34300
rect 9355 34244 9411 34300
rect 9411 34244 9415 34300
rect 9351 34240 9415 34244
rect 3004 33764 3068 33828
rect 4215 33756 4279 33760
rect 4215 33700 4219 33756
rect 4219 33700 4275 33756
rect 4275 33700 4279 33756
rect 4215 33696 4279 33700
rect 4295 33756 4359 33760
rect 4295 33700 4299 33756
rect 4299 33700 4355 33756
rect 4355 33700 4359 33756
rect 4295 33696 4359 33700
rect 4375 33756 4439 33760
rect 4375 33700 4379 33756
rect 4379 33700 4435 33756
rect 4435 33700 4439 33756
rect 4375 33696 4439 33700
rect 4455 33756 4519 33760
rect 4455 33700 4459 33756
rect 4459 33700 4515 33756
rect 4515 33700 4519 33756
rect 4455 33696 4519 33700
rect 7479 33756 7543 33760
rect 7479 33700 7483 33756
rect 7483 33700 7539 33756
rect 7539 33700 7543 33756
rect 7479 33696 7543 33700
rect 7559 33756 7623 33760
rect 7559 33700 7563 33756
rect 7563 33700 7619 33756
rect 7619 33700 7623 33756
rect 7559 33696 7623 33700
rect 7639 33756 7703 33760
rect 7639 33700 7643 33756
rect 7643 33700 7699 33756
rect 7699 33700 7703 33756
rect 7639 33696 7703 33700
rect 7719 33756 7783 33760
rect 7719 33700 7723 33756
rect 7723 33700 7779 33756
rect 7779 33700 7783 33756
rect 7719 33696 7783 33700
rect 2584 33212 2648 33216
rect 2584 33156 2588 33212
rect 2588 33156 2644 33212
rect 2644 33156 2648 33212
rect 2584 33152 2648 33156
rect 2664 33212 2728 33216
rect 2664 33156 2668 33212
rect 2668 33156 2724 33212
rect 2724 33156 2728 33212
rect 2664 33152 2728 33156
rect 2744 33212 2808 33216
rect 2744 33156 2748 33212
rect 2748 33156 2804 33212
rect 2804 33156 2808 33212
rect 2744 33152 2808 33156
rect 2824 33212 2888 33216
rect 2824 33156 2828 33212
rect 2828 33156 2884 33212
rect 2884 33156 2888 33212
rect 2824 33152 2888 33156
rect 5847 33212 5911 33216
rect 5847 33156 5851 33212
rect 5851 33156 5907 33212
rect 5907 33156 5911 33212
rect 5847 33152 5911 33156
rect 5927 33212 5991 33216
rect 5927 33156 5931 33212
rect 5931 33156 5987 33212
rect 5987 33156 5991 33212
rect 5927 33152 5991 33156
rect 6007 33212 6071 33216
rect 6007 33156 6011 33212
rect 6011 33156 6067 33212
rect 6067 33156 6071 33212
rect 6007 33152 6071 33156
rect 6087 33212 6151 33216
rect 6087 33156 6091 33212
rect 6091 33156 6147 33212
rect 6147 33156 6151 33212
rect 6087 33152 6151 33156
rect 9111 33212 9175 33216
rect 9111 33156 9115 33212
rect 9115 33156 9171 33212
rect 9171 33156 9175 33212
rect 9111 33152 9175 33156
rect 9191 33212 9255 33216
rect 9191 33156 9195 33212
rect 9195 33156 9251 33212
rect 9251 33156 9255 33212
rect 9191 33152 9255 33156
rect 9271 33212 9335 33216
rect 9271 33156 9275 33212
rect 9275 33156 9331 33212
rect 9331 33156 9335 33212
rect 9271 33152 9335 33156
rect 9351 33212 9415 33216
rect 9351 33156 9355 33212
rect 9355 33156 9411 33212
rect 9411 33156 9415 33212
rect 9351 33152 9415 33156
rect 4215 32668 4279 32672
rect 4215 32612 4219 32668
rect 4219 32612 4275 32668
rect 4275 32612 4279 32668
rect 4215 32608 4279 32612
rect 4295 32668 4359 32672
rect 4295 32612 4299 32668
rect 4299 32612 4355 32668
rect 4355 32612 4359 32668
rect 4295 32608 4359 32612
rect 4375 32668 4439 32672
rect 4375 32612 4379 32668
rect 4379 32612 4435 32668
rect 4435 32612 4439 32668
rect 4375 32608 4439 32612
rect 4455 32668 4519 32672
rect 4455 32612 4459 32668
rect 4459 32612 4515 32668
rect 4515 32612 4519 32668
rect 4455 32608 4519 32612
rect 7479 32668 7543 32672
rect 7479 32612 7483 32668
rect 7483 32612 7539 32668
rect 7539 32612 7543 32668
rect 7479 32608 7543 32612
rect 7559 32668 7623 32672
rect 7559 32612 7563 32668
rect 7563 32612 7619 32668
rect 7619 32612 7623 32668
rect 7559 32608 7623 32612
rect 7639 32668 7703 32672
rect 7639 32612 7643 32668
rect 7643 32612 7699 32668
rect 7699 32612 7703 32668
rect 7639 32608 7703 32612
rect 7719 32668 7783 32672
rect 7719 32612 7723 32668
rect 7723 32612 7779 32668
rect 7779 32612 7783 32668
rect 7719 32608 7783 32612
rect 2268 32600 2332 32604
rect 2268 32544 2318 32600
rect 2318 32544 2332 32600
rect 2268 32540 2332 32544
rect 2084 32404 2148 32468
rect 2584 32124 2648 32128
rect 2584 32068 2588 32124
rect 2588 32068 2644 32124
rect 2644 32068 2648 32124
rect 2584 32064 2648 32068
rect 2664 32124 2728 32128
rect 2664 32068 2668 32124
rect 2668 32068 2724 32124
rect 2724 32068 2728 32124
rect 2664 32064 2728 32068
rect 2744 32124 2808 32128
rect 2744 32068 2748 32124
rect 2748 32068 2804 32124
rect 2804 32068 2808 32124
rect 2744 32064 2808 32068
rect 2824 32124 2888 32128
rect 2824 32068 2828 32124
rect 2828 32068 2884 32124
rect 2884 32068 2888 32124
rect 2824 32064 2888 32068
rect 5847 32124 5911 32128
rect 5847 32068 5851 32124
rect 5851 32068 5907 32124
rect 5907 32068 5911 32124
rect 5847 32064 5911 32068
rect 5927 32124 5991 32128
rect 5927 32068 5931 32124
rect 5931 32068 5987 32124
rect 5987 32068 5991 32124
rect 5927 32064 5991 32068
rect 6007 32124 6071 32128
rect 6007 32068 6011 32124
rect 6011 32068 6067 32124
rect 6067 32068 6071 32124
rect 6007 32064 6071 32068
rect 6087 32124 6151 32128
rect 6087 32068 6091 32124
rect 6091 32068 6147 32124
rect 6147 32068 6151 32124
rect 6087 32064 6151 32068
rect 9111 32124 9175 32128
rect 9111 32068 9115 32124
rect 9115 32068 9171 32124
rect 9171 32068 9175 32124
rect 9111 32064 9175 32068
rect 9191 32124 9255 32128
rect 9191 32068 9195 32124
rect 9195 32068 9251 32124
rect 9251 32068 9255 32124
rect 9191 32064 9255 32068
rect 9271 32124 9335 32128
rect 9271 32068 9275 32124
rect 9275 32068 9331 32124
rect 9331 32068 9335 32124
rect 9271 32064 9335 32068
rect 9351 32124 9415 32128
rect 9351 32068 9355 32124
rect 9355 32068 9411 32124
rect 9411 32068 9415 32124
rect 9351 32064 9415 32068
rect 1532 31996 1596 32060
rect 1716 31784 1780 31788
rect 1716 31728 1766 31784
rect 1766 31728 1780 31784
rect 1716 31724 1780 31728
rect 3556 31648 3620 31652
rect 3556 31592 3606 31648
rect 3606 31592 3620 31648
rect 3556 31588 3620 31592
rect 4215 31580 4279 31584
rect 4215 31524 4219 31580
rect 4219 31524 4275 31580
rect 4275 31524 4279 31580
rect 4215 31520 4279 31524
rect 4295 31580 4359 31584
rect 4295 31524 4299 31580
rect 4299 31524 4355 31580
rect 4355 31524 4359 31580
rect 4295 31520 4359 31524
rect 4375 31580 4439 31584
rect 4375 31524 4379 31580
rect 4379 31524 4435 31580
rect 4435 31524 4439 31580
rect 4375 31520 4439 31524
rect 4455 31580 4519 31584
rect 4455 31524 4459 31580
rect 4459 31524 4515 31580
rect 4515 31524 4519 31580
rect 4455 31520 4519 31524
rect 7479 31580 7543 31584
rect 7479 31524 7483 31580
rect 7483 31524 7539 31580
rect 7539 31524 7543 31580
rect 7479 31520 7543 31524
rect 7559 31580 7623 31584
rect 7559 31524 7563 31580
rect 7563 31524 7619 31580
rect 7619 31524 7623 31580
rect 7559 31520 7623 31524
rect 7639 31580 7703 31584
rect 7639 31524 7643 31580
rect 7643 31524 7699 31580
rect 7699 31524 7703 31580
rect 7639 31520 7703 31524
rect 7719 31580 7783 31584
rect 7719 31524 7723 31580
rect 7723 31524 7779 31580
rect 7779 31524 7783 31580
rect 7719 31520 7783 31524
rect 2584 31036 2648 31040
rect 2584 30980 2588 31036
rect 2588 30980 2644 31036
rect 2644 30980 2648 31036
rect 2584 30976 2648 30980
rect 2664 31036 2728 31040
rect 2664 30980 2668 31036
rect 2668 30980 2724 31036
rect 2724 30980 2728 31036
rect 2664 30976 2728 30980
rect 2744 31036 2808 31040
rect 2744 30980 2748 31036
rect 2748 30980 2804 31036
rect 2804 30980 2808 31036
rect 2744 30976 2808 30980
rect 2824 31036 2888 31040
rect 2824 30980 2828 31036
rect 2828 30980 2884 31036
rect 2884 30980 2888 31036
rect 2824 30976 2888 30980
rect 5847 31036 5911 31040
rect 5847 30980 5851 31036
rect 5851 30980 5907 31036
rect 5907 30980 5911 31036
rect 5847 30976 5911 30980
rect 5927 31036 5991 31040
rect 5927 30980 5931 31036
rect 5931 30980 5987 31036
rect 5987 30980 5991 31036
rect 5927 30976 5991 30980
rect 6007 31036 6071 31040
rect 6007 30980 6011 31036
rect 6011 30980 6067 31036
rect 6067 30980 6071 31036
rect 6007 30976 6071 30980
rect 6087 31036 6151 31040
rect 6087 30980 6091 31036
rect 6091 30980 6147 31036
rect 6147 30980 6151 31036
rect 6087 30976 6151 30980
rect 9111 31036 9175 31040
rect 9111 30980 9115 31036
rect 9115 30980 9171 31036
rect 9171 30980 9175 31036
rect 9111 30976 9175 30980
rect 9191 31036 9255 31040
rect 9191 30980 9195 31036
rect 9195 30980 9251 31036
rect 9251 30980 9255 31036
rect 9191 30976 9255 30980
rect 9271 31036 9335 31040
rect 9271 30980 9275 31036
rect 9275 30980 9331 31036
rect 9331 30980 9335 31036
rect 9271 30976 9335 30980
rect 9351 31036 9415 31040
rect 9351 30980 9355 31036
rect 9355 30980 9411 31036
rect 9411 30980 9415 31036
rect 9351 30976 9415 30980
rect 4215 30492 4279 30496
rect 4215 30436 4219 30492
rect 4219 30436 4275 30492
rect 4275 30436 4279 30492
rect 4215 30432 4279 30436
rect 4295 30492 4359 30496
rect 4295 30436 4299 30492
rect 4299 30436 4355 30492
rect 4355 30436 4359 30492
rect 4295 30432 4359 30436
rect 4375 30492 4439 30496
rect 4375 30436 4379 30492
rect 4379 30436 4435 30492
rect 4435 30436 4439 30492
rect 4375 30432 4439 30436
rect 4455 30492 4519 30496
rect 4455 30436 4459 30492
rect 4459 30436 4515 30492
rect 4515 30436 4519 30492
rect 4455 30432 4519 30436
rect 7479 30492 7543 30496
rect 7479 30436 7483 30492
rect 7483 30436 7539 30492
rect 7539 30436 7543 30492
rect 7479 30432 7543 30436
rect 7559 30492 7623 30496
rect 7559 30436 7563 30492
rect 7563 30436 7619 30492
rect 7619 30436 7623 30492
rect 7559 30432 7623 30436
rect 7639 30492 7703 30496
rect 7639 30436 7643 30492
rect 7643 30436 7699 30492
rect 7699 30436 7703 30492
rect 7639 30432 7703 30436
rect 7719 30492 7783 30496
rect 7719 30436 7723 30492
rect 7723 30436 7779 30492
rect 7779 30436 7783 30492
rect 7719 30432 7783 30436
rect 2584 29948 2648 29952
rect 2584 29892 2588 29948
rect 2588 29892 2644 29948
rect 2644 29892 2648 29948
rect 2584 29888 2648 29892
rect 2664 29948 2728 29952
rect 2664 29892 2668 29948
rect 2668 29892 2724 29948
rect 2724 29892 2728 29948
rect 2664 29888 2728 29892
rect 2744 29948 2808 29952
rect 2744 29892 2748 29948
rect 2748 29892 2804 29948
rect 2804 29892 2808 29948
rect 2744 29888 2808 29892
rect 2824 29948 2888 29952
rect 2824 29892 2828 29948
rect 2828 29892 2884 29948
rect 2884 29892 2888 29948
rect 2824 29888 2888 29892
rect 5847 29948 5911 29952
rect 5847 29892 5851 29948
rect 5851 29892 5907 29948
rect 5907 29892 5911 29948
rect 5847 29888 5911 29892
rect 5927 29948 5991 29952
rect 5927 29892 5931 29948
rect 5931 29892 5987 29948
rect 5987 29892 5991 29948
rect 5927 29888 5991 29892
rect 6007 29948 6071 29952
rect 6007 29892 6011 29948
rect 6011 29892 6067 29948
rect 6067 29892 6071 29948
rect 6007 29888 6071 29892
rect 6087 29948 6151 29952
rect 6087 29892 6091 29948
rect 6091 29892 6147 29948
rect 6147 29892 6151 29948
rect 6087 29888 6151 29892
rect 9111 29948 9175 29952
rect 9111 29892 9115 29948
rect 9115 29892 9171 29948
rect 9171 29892 9175 29948
rect 9111 29888 9175 29892
rect 9191 29948 9255 29952
rect 9191 29892 9195 29948
rect 9195 29892 9251 29948
rect 9251 29892 9255 29948
rect 9191 29888 9255 29892
rect 9271 29948 9335 29952
rect 9271 29892 9275 29948
rect 9275 29892 9331 29948
rect 9331 29892 9335 29948
rect 9271 29888 9335 29892
rect 9351 29948 9415 29952
rect 9351 29892 9355 29948
rect 9355 29892 9411 29948
rect 9411 29892 9415 29948
rect 9351 29888 9415 29892
rect 4215 29404 4279 29408
rect 4215 29348 4219 29404
rect 4219 29348 4275 29404
rect 4275 29348 4279 29404
rect 4215 29344 4279 29348
rect 4295 29404 4359 29408
rect 4295 29348 4299 29404
rect 4299 29348 4355 29404
rect 4355 29348 4359 29404
rect 4295 29344 4359 29348
rect 4375 29404 4439 29408
rect 4375 29348 4379 29404
rect 4379 29348 4435 29404
rect 4435 29348 4439 29404
rect 4375 29344 4439 29348
rect 4455 29404 4519 29408
rect 4455 29348 4459 29404
rect 4459 29348 4515 29404
rect 4515 29348 4519 29404
rect 4455 29344 4519 29348
rect 7479 29404 7543 29408
rect 7479 29348 7483 29404
rect 7483 29348 7539 29404
rect 7539 29348 7543 29404
rect 7479 29344 7543 29348
rect 7559 29404 7623 29408
rect 7559 29348 7563 29404
rect 7563 29348 7619 29404
rect 7619 29348 7623 29404
rect 7559 29344 7623 29348
rect 7639 29404 7703 29408
rect 7639 29348 7643 29404
rect 7643 29348 7699 29404
rect 7699 29348 7703 29404
rect 7639 29344 7703 29348
rect 7719 29404 7783 29408
rect 7719 29348 7723 29404
rect 7723 29348 7779 29404
rect 7779 29348 7783 29404
rect 7719 29344 7783 29348
rect 1716 29200 1780 29204
rect 1716 29144 1766 29200
rect 1766 29144 1780 29200
rect 1716 29140 1780 29144
rect 3004 28868 3068 28932
rect 2584 28860 2648 28864
rect 2584 28804 2588 28860
rect 2588 28804 2644 28860
rect 2644 28804 2648 28860
rect 2584 28800 2648 28804
rect 2664 28860 2728 28864
rect 2664 28804 2668 28860
rect 2668 28804 2724 28860
rect 2724 28804 2728 28860
rect 2664 28800 2728 28804
rect 2744 28860 2808 28864
rect 2744 28804 2748 28860
rect 2748 28804 2804 28860
rect 2804 28804 2808 28860
rect 2744 28800 2808 28804
rect 2824 28860 2888 28864
rect 2824 28804 2828 28860
rect 2828 28804 2884 28860
rect 2884 28804 2888 28860
rect 2824 28800 2888 28804
rect 5847 28860 5911 28864
rect 5847 28804 5851 28860
rect 5851 28804 5907 28860
rect 5907 28804 5911 28860
rect 5847 28800 5911 28804
rect 5927 28860 5991 28864
rect 5927 28804 5931 28860
rect 5931 28804 5987 28860
rect 5987 28804 5991 28860
rect 5927 28800 5991 28804
rect 6007 28860 6071 28864
rect 6007 28804 6011 28860
rect 6011 28804 6067 28860
rect 6067 28804 6071 28860
rect 6007 28800 6071 28804
rect 6087 28860 6151 28864
rect 6087 28804 6091 28860
rect 6091 28804 6147 28860
rect 6147 28804 6151 28860
rect 6087 28800 6151 28804
rect 9111 28860 9175 28864
rect 9111 28804 9115 28860
rect 9115 28804 9171 28860
rect 9171 28804 9175 28860
rect 9111 28800 9175 28804
rect 9191 28860 9255 28864
rect 9191 28804 9195 28860
rect 9195 28804 9251 28860
rect 9251 28804 9255 28860
rect 9191 28800 9255 28804
rect 9271 28860 9335 28864
rect 9271 28804 9275 28860
rect 9275 28804 9331 28860
rect 9331 28804 9335 28860
rect 9271 28800 9335 28804
rect 9351 28860 9415 28864
rect 9351 28804 9355 28860
rect 9355 28804 9411 28860
rect 9411 28804 9415 28860
rect 9351 28800 9415 28804
rect 4215 28316 4279 28320
rect 4215 28260 4219 28316
rect 4219 28260 4275 28316
rect 4275 28260 4279 28316
rect 4215 28256 4279 28260
rect 4295 28316 4359 28320
rect 4295 28260 4299 28316
rect 4299 28260 4355 28316
rect 4355 28260 4359 28316
rect 4295 28256 4359 28260
rect 4375 28316 4439 28320
rect 4375 28260 4379 28316
rect 4379 28260 4435 28316
rect 4435 28260 4439 28316
rect 4375 28256 4439 28260
rect 4455 28316 4519 28320
rect 4455 28260 4459 28316
rect 4459 28260 4515 28316
rect 4515 28260 4519 28316
rect 4455 28256 4519 28260
rect 7479 28316 7543 28320
rect 7479 28260 7483 28316
rect 7483 28260 7539 28316
rect 7539 28260 7543 28316
rect 7479 28256 7543 28260
rect 7559 28316 7623 28320
rect 7559 28260 7563 28316
rect 7563 28260 7619 28316
rect 7619 28260 7623 28316
rect 7559 28256 7623 28260
rect 7639 28316 7703 28320
rect 7639 28260 7643 28316
rect 7643 28260 7699 28316
rect 7699 28260 7703 28316
rect 7639 28256 7703 28260
rect 7719 28316 7783 28320
rect 7719 28260 7723 28316
rect 7723 28260 7779 28316
rect 7779 28260 7783 28316
rect 7719 28256 7783 28260
rect 2584 27772 2648 27776
rect 2584 27716 2588 27772
rect 2588 27716 2644 27772
rect 2644 27716 2648 27772
rect 2584 27712 2648 27716
rect 2664 27772 2728 27776
rect 2664 27716 2668 27772
rect 2668 27716 2724 27772
rect 2724 27716 2728 27772
rect 2664 27712 2728 27716
rect 2744 27772 2808 27776
rect 2744 27716 2748 27772
rect 2748 27716 2804 27772
rect 2804 27716 2808 27772
rect 2744 27712 2808 27716
rect 2824 27772 2888 27776
rect 2824 27716 2828 27772
rect 2828 27716 2884 27772
rect 2884 27716 2888 27772
rect 2824 27712 2888 27716
rect 5847 27772 5911 27776
rect 5847 27716 5851 27772
rect 5851 27716 5907 27772
rect 5907 27716 5911 27772
rect 5847 27712 5911 27716
rect 5927 27772 5991 27776
rect 5927 27716 5931 27772
rect 5931 27716 5987 27772
rect 5987 27716 5991 27772
rect 5927 27712 5991 27716
rect 6007 27772 6071 27776
rect 6007 27716 6011 27772
rect 6011 27716 6067 27772
rect 6067 27716 6071 27772
rect 6007 27712 6071 27716
rect 6087 27772 6151 27776
rect 6087 27716 6091 27772
rect 6091 27716 6147 27772
rect 6147 27716 6151 27772
rect 6087 27712 6151 27716
rect 9111 27772 9175 27776
rect 9111 27716 9115 27772
rect 9115 27716 9171 27772
rect 9171 27716 9175 27772
rect 9111 27712 9175 27716
rect 9191 27772 9255 27776
rect 9191 27716 9195 27772
rect 9195 27716 9251 27772
rect 9251 27716 9255 27772
rect 9191 27712 9255 27716
rect 9271 27772 9335 27776
rect 9271 27716 9275 27772
rect 9275 27716 9331 27772
rect 9331 27716 9335 27772
rect 9271 27712 9335 27716
rect 9351 27772 9415 27776
rect 9351 27716 9355 27772
rect 9355 27716 9411 27772
rect 9411 27716 9415 27772
rect 9351 27712 9415 27716
rect 4215 27228 4279 27232
rect 4215 27172 4219 27228
rect 4219 27172 4275 27228
rect 4275 27172 4279 27228
rect 4215 27168 4279 27172
rect 4295 27228 4359 27232
rect 4295 27172 4299 27228
rect 4299 27172 4355 27228
rect 4355 27172 4359 27228
rect 4295 27168 4359 27172
rect 4375 27228 4439 27232
rect 4375 27172 4379 27228
rect 4379 27172 4435 27228
rect 4435 27172 4439 27228
rect 4375 27168 4439 27172
rect 4455 27228 4519 27232
rect 4455 27172 4459 27228
rect 4459 27172 4515 27228
rect 4515 27172 4519 27228
rect 4455 27168 4519 27172
rect 7479 27228 7543 27232
rect 7479 27172 7483 27228
rect 7483 27172 7539 27228
rect 7539 27172 7543 27228
rect 7479 27168 7543 27172
rect 7559 27228 7623 27232
rect 7559 27172 7563 27228
rect 7563 27172 7619 27228
rect 7619 27172 7623 27228
rect 7559 27168 7623 27172
rect 7639 27228 7703 27232
rect 7639 27172 7643 27228
rect 7643 27172 7699 27228
rect 7699 27172 7703 27228
rect 7639 27168 7703 27172
rect 7719 27228 7783 27232
rect 7719 27172 7723 27228
rect 7723 27172 7779 27228
rect 7779 27172 7783 27228
rect 7719 27168 7783 27172
rect 3004 26692 3068 26756
rect 2584 26684 2648 26688
rect 2584 26628 2588 26684
rect 2588 26628 2644 26684
rect 2644 26628 2648 26684
rect 2584 26624 2648 26628
rect 2664 26684 2728 26688
rect 2664 26628 2668 26684
rect 2668 26628 2724 26684
rect 2724 26628 2728 26684
rect 2664 26624 2728 26628
rect 2744 26684 2808 26688
rect 2744 26628 2748 26684
rect 2748 26628 2804 26684
rect 2804 26628 2808 26684
rect 2744 26624 2808 26628
rect 2824 26684 2888 26688
rect 2824 26628 2828 26684
rect 2828 26628 2884 26684
rect 2884 26628 2888 26684
rect 2824 26624 2888 26628
rect 5847 26684 5911 26688
rect 5847 26628 5851 26684
rect 5851 26628 5907 26684
rect 5907 26628 5911 26684
rect 5847 26624 5911 26628
rect 5927 26684 5991 26688
rect 5927 26628 5931 26684
rect 5931 26628 5987 26684
rect 5987 26628 5991 26684
rect 5927 26624 5991 26628
rect 6007 26684 6071 26688
rect 6007 26628 6011 26684
rect 6011 26628 6067 26684
rect 6067 26628 6071 26684
rect 6007 26624 6071 26628
rect 6087 26684 6151 26688
rect 6087 26628 6091 26684
rect 6091 26628 6147 26684
rect 6147 26628 6151 26684
rect 6087 26624 6151 26628
rect 9111 26684 9175 26688
rect 9111 26628 9115 26684
rect 9115 26628 9171 26684
rect 9171 26628 9175 26684
rect 9111 26624 9175 26628
rect 9191 26684 9255 26688
rect 9191 26628 9195 26684
rect 9195 26628 9251 26684
rect 9251 26628 9255 26684
rect 9191 26624 9255 26628
rect 9271 26684 9335 26688
rect 9271 26628 9275 26684
rect 9275 26628 9331 26684
rect 9331 26628 9335 26684
rect 9271 26624 9335 26628
rect 9351 26684 9415 26688
rect 9351 26628 9355 26684
rect 9355 26628 9411 26684
rect 9411 26628 9415 26684
rect 9351 26624 9415 26628
rect 4215 26140 4279 26144
rect 4215 26084 4219 26140
rect 4219 26084 4275 26140
rect 4275 26084 4279 26140
rect 4215 26080 4279 26084
rect 4295 26140 4359 26144
rect 4295 26084 4299 26140
rect 4299 26084 4355 26140
rect 4355 26084 4359 26140
rect 4295 26080 4359 26084
rect 4375 26140 4439 26144
rect 4375 26084 4379 26140
rect 4379 26084 4435 26140
rect 4435 26084 4439 26140
rect 4375 26080 4439 26084
rect 4455 26140 4519 26144
rect 4455 26084 4459 26140
rect 4459 26084 4515 26140
rect 4515 26084 4519 26140
rect 4455 26080 4519 26084
rect 7479 26140 7543 26144
rect 7479 26084 7483 26140
rect 7483 26084 7539 26140
rect 7539 26084 7543 26140
rect 7479 26080 7543 26084
rect 7559 26140 7623 26144
rect 7559 26084 7563 26140
rect 7563 26084 7619 26140
rect 7619 26084 7623 26140
rect 7559 26080 7623 26084
rect 7639 26140 7703 26144
rect 7639 26084 7643 26140
rect 7643 26084 7699 26140
rect 7699 26084 7703 26140
rect 7639 26080 7703 26084
rect 7719 26140 7783 26144
rect 7719 26084 7723 26140
rect 7723 26084 7779 26140
rect 7779 26084 7783 26140
rect 7719 26080 7783 26084
rect 2584 25596 2648 25600
rect 2584 25540 2588 25596
rect 2588 25540 2644 25596
rect 2644 25540 2648 25596
rect 2584 25536 2648 25540
rect 2664 25596 2728 25600
rect 2664 25540 2668 25596
rect 2668 25540 2724 25596
rect 2724 25540 2728 25596
rect 2664 25536 2728 25540
rect 2744 25596 2808 25600
rect 2744 25540 2748 25596
rect 2748 25540 2804 25596
rect 2804 25540 2808 25596
rect 2744 25536 2808 25540
rect 2824 25596 2888 25600
rect 2824 25540 2828 25596
rect 2828 25540 2884 25596
rect 2884 25540 2888 25596
rect 2824 25536 2888 25540
rect 5847 25596 5911 25600
rect 5847 25540 5851 25596
rect 5851 25540 5907 25596
rect 5907 25540 5911 25596
rect 5847 25536 5911 25540
rect 5927 25596 5991 25600
rect 5927 25540 5931 25596
rect 5931 25540 5987 25596
rect 5987 25540 5991 25596
rect 5927 25536 5991 25540
rect 6007 25596 6071 25600
rect 6007 25540 6011 25596
rect 6011 25540 6067 25596
rect 6067 25540 6071 25596
rect 6007 25536 6071 25540
rect 6087 25596 6151 25600
rect 6087 25540 6091 25596
rect 6091 25540 6147 25596
rect 6147 25540 6151 25596
rect 6087 25536 6151 25540
rect 9111 25596 9175 25600
rect 9111 25540 9115 25596
rect 9115 25540 9171 25596
rect 9171 25540 9175 25596
rect 9111 25536 9175 25540
rect 9191 25596 9255 25600
rect 9191 25540 9195 25596
rect 9195 25540 9251 25596
rect 9251 25540 9255 25596
rect 9191 25536 9255 25540
rect 9271 25596 9335 25600
rect 9271 25540 9275 25596
rect 9275 25540 9331 25596
rect 9331 25540 9335 25596
rect 9271 25536 9335 25540
rect 9351 25596 9415 25600
rect 9351 25540 9355 25596
rect 9355 25540 9411 25596
rect 9411 25540 9415 25596
rect 9351 25536 9415 25540
rect 4215 25052 4279 25056
rect 4215 24996 4219 25052
rect 4219 24996 4275 25052
rect 4275 24996 4279 25052
rect 4215 24992 4279 24996
rect 4295 25052 4359 25056
rect 4295 24996 4299 25052
rect 4299 24996 4355 25052
rect 4355 24996 4359 25052
rect 4295 24992 4359 24996
rect 4375 25052 4439 25056
rect 4375 24996 4379 25052
rect 4379 24996 4435 25052
rect 4435 24996 4439 25052
rect 4375 24992 4439 24996
rect 4455 25052 4519 25056
rect 4455 24996 4459 25052
rect 4459 24996 4515 25052
rect 4515 24996 4519 25052
rect 4455 24992 4519 24996
rect 7479 25052 7543 25056
rect 7479 24996 7483 25052
rect 7483 24996 7539 25052
rect 7539 24996 7543 25052
rect 7479 24992 7543 24996
rect 7559 25052 7623 25056
rect 7559 24996 7563 25052
rect 7563 24996 7619 25052
rect 7619 24996 7623 25052
rect 7559 24992 7623 24996
rect 7639 25052 7703 25056
rect 7639 24996 7643 25052
rect 7643 24996 7699 25052
rect 7699 24996 7703 25052
rect 7639 24992 7703 24996
rect 7719 25052 7783 25056
rect 7719 24996 7723 25052
rect 7723 24996 7779 25052
rect 7779 24996 7783 25052
rect 7719 24992 7783 24996
rect 2584 24508 2648 24512
rect 2584 24452 2588 24508
rect 2588 24452 2644 24508
rect 2644 24452 2648 24508
rect 2584 24448 2648 24452
rect 2664 24508 2728 24512
rect 2664 24452 2668 24508
rect 2668 24452 2724 24508
rect 2724 24452 2728 24508
rect 2664 24448 2728 24452
rect 2744 24508 2808 24512
rect 2744 24452 2748 24508
rect 2748 24452 2804 24508
rect 2804 24452 2808 24508
rect 2744 24448 2808 24452
rect 2824 24508 2888 24512
rect 2824 24452 2828 24508
rect 2828 24452 2884 24508
rect 2884 24452 2888 24508
rect 2824 24448 2888 24452
rect 5847 24508 5911 24512
rect 5847 24452 5851 24508
rect 5851 24452 5907 24508
rect 5907 24452 5911 24508
rect 5847 24448 5911 24452
rect 5927 24508 5991 24512
rect 5927 24452 5931 24508
rect 5931 24452 5987 24508
rect 5987 24452 5991 24508
rect 5927 24448 5991 24452
rect 6007 24508 6071 24512
rect 6007 24452 6011 24508
rect 6011 24452 6067 24508
rect 6067 24452 6071 24508
rect 6007 24448 6071 24452
rect 6087 24508 6151 24512
rect 6087 24452 6091 24508
rect 6091 24452 6147 24508
rect 6147 24452 6151 24508
rect 6087 24448 6151 24452
rect 9111 24508 9175 24512
rect 9111 24452 9115 24508
rect 9115 24452 9171 24508
rect 9171 24452 9175 24508
rect 9111 24448 9175 24452
rect 9191 24508 9255 24512
rect 9191 24452 9195 24508
rect 9195 24452 9251 24508
rect 9251 24452 9255 24508
rect 9191 24448 9255 24452
rect 9271 24508 9335 24512
rect 9271 24452 9275 24508
rect 9275 24452 9331 24508
rect 9331 24452 9335 24508
rect 9271 24448 9335 24452
rect 9351 24508 9415 24512
rect 9351 24452 9355 24508
rect 9355 24452 9411 24508
rect 9411 24452 9415 24508
rect 9351 24448 9415 24452
rect 4215 23964 4279 23968
rect 4215 23908 4219 23964
rect 4219 23908 4275 23964
rect 4275 23908 4279 23964
rect 4215 23904 4279 23908
rect 4295 23964 4359 23968
rect 4295 23908 4299 23964
rect 4299 23908 4355 23964
rect 4355 23908 4359 23964
rect 4295 23904 4359 23908
rect 4375 23964 4439 23968
rect 4375 23908 4379 23964
rect 4379 23908 4435 23964
rect 4435 23908 4439 23964
rect 4375 23904 4439 23908
rect 4455 23964 4519 23968
rect 4455 23908 4459 23964
rect 4459 23908 4515 23964
rect 4515 23908 4519 23964
rect 4455 23904 4519 23908
rect 7479 23964 7543 23968
rect 7479 23908 7483 23964
rect 7483 23908 7539 23964
rect 7539 23908 7543 23964
rect 7479 23904 7543 23908
rect 7559 23964 7623 23968
rect 7559 23908 7563 23964
rect 7563 23908 7619 23964
rect 7619 23908 7623 23964
rect 7559 23904 7623 23908
rect 7639 23964 7703 23968
rect 7639 23908 7643 23964
rect 7643 23908 7699 23964
rect 7699 23908 7703 23964
rect 7639 23904 7703 23908
rect 7719 23964 7783 23968
rect 7719 23908 7723 23964
rect 7723 23908 7779 23964
rect 7779 23908 7783 23964
rect 7719 23904 7783 23908
rect 2584 23420 2648 23424
rect 2584 23364 2588 23420
rect 2588 23364 2644 23420
rect 2644 23364 2648 23420
rect 2584 23360 2648 23364
rect 2664 23420 2728 23424
rect 2664 23364 2668 23420
rect 2668 23364 2724 23420
rect 2724 23364 2728 23420
rect 2664 23360 2728 23364
rect 2744 23420 2808 23424
rect 2744 23364 2748 23420
rect 2748 23364 2804 23420
rect 2804 23364 2808 23420
rect 2744 23360 2808 23364
rect 2824 23420 2888 23424
rect 2824 23364 2828 23420
rect 2828 23364 2884 23420
rect 2884 23364 2888 23420
rect 2824 23360 2888 23364
rect 5847 23420 5911 23424
rect 5847 23364 5851 23420
rect 5851 23364 5907 23420
rect 5907 23364 5911 23420
rect 5847 23360 5911 23364
rect 5927 23420 5991 23424
rect 5927 23364 5931 23420
rect 5931 23364 5987 23420
rect 5987 23364 5991 23420
rect 5927 23360 5991 23364
rect 6007 23420 6071 23424
rect 6007 23364 6011 23420
rect 6011 23364 6067 23420
rect 6067 23364 6071 23420
rect 6007 23360 6071 23364
rect 6087 23420 6151 23424
rect 6087 23364 6091 23420
rect 6091 23364 6147 23420
rect 6147 23364 6151 23420
rect 6087 23360 6151 23364
rect 9111 23420 9175 23424
rect 9111 23364 9115 23420
rect 9115 23364 9171 23420
rect 9171 23364 9175 23420
rect 9111 23360 9175 23364
rect 9191 23420 9255 23424
rect 9191 23364 9195 23420
rect 9195 23364 9251 23420
rect 9251 23364 9255 23420
rect 9191 23360 9255 23364
rect 9271 23420 9335 23424
rect 9271 23364 9275 23420
rect 9275 23364 9331 23420
rect 9331 23364 9335 23420
rect 9271 23360 9335 23364
rect 9351 23420 9415 23424
rect 9351 23364 9355 23420
rect 9355 23364 9411 23420
rect 9411 23364 9415 23420
rect 9351 23360 9415 23364
rect 4215 22876 4279 22880
rect 4215 22820 4219 22876
rect 4219 22820 4275 22876
rect 4275 22820 4279 22876
rect 4215 22816 4279 22820
rect 4295 22876 4359 22880
rect 4295 22820 4299 22876
rect 4299 22820 4355 22876
rect 4355 22820 4359 22876
rect 4295 22816 4359 22820
rect 4375 22876 4439 22880
rect 4375 22820 4379 22876
rect 4379 22820 4435 22876
rect 4435 22820 4439 22876
rect 4375 22816 4439 22820
rect 4455 22876 4519 22880
rect 4455 22820 4459 22876
rect 4459 22820 4515 22876
rect 4515 22820 4519 22876
rect 4455 22816 4519 22820
rect 7479 22876 7543 22880
rect 7479 22820 7483 22876
rect 7483 22820 7539 22876
rect 7539 22820 7543 22876
rect 7479 22816 7543 22820
rect 7559 22876 7623 22880
rect 7559 22820 7563 22876
rect 7563 22820 7619 22876
rect 7619 22820 7623 22876
rect 7559 22816 7623 22820
rect 7639 22876 7703 22880
rect 7639 22820 7643 22876
rect 7643 22820 7699 22876
rect 7699 22820 7703 22876
rect 7639 22816 7703 22820
rect 7719 22876 7783 22880
rect 7719 22820 7723 22876
rect 7723 22820 7779 22876
rect 7779 22820 7783 22876
rect 7719 22816 7783 22820
rect 2584 22332 2648 22336
rect 2584 22276 2588 22332
rect 2588 22276 2644 22332
rect 2644 22276 2648 22332
rect 2584 22272 2648 22276
rect 2664 22332 2728 22336
rect 2664 22276 2668 22332
rect 2668 22276 2724 22332
rect 2724 22276 2728 22332
rect 2664 22272 2728 22276
rect 2744 22332 2808 22336
rect 2744 22276 2748 22332
rect 2748 22276 2804 22332
rect 2804 22276 2808 22332
rect 2744 22272 2808 22276
rect 2824 22332 2888 22336
rect 2824 22276 2828 22332
rect 2828 22276 2884 22332
rect 2884 22276 2888 22332
rect 2824 22272 2888 22276
rect 5847 22332 5911 22336
rect 5847 22276 5851 22332
rect 5851 22276 5907 22332
rect 5907 22276 5911 22332
rect 5847 22272 5911 22276
rect 5927 22332 5991 22336
rect 5927 22276 5931 22332
rect 5931 22276 5987 22332
rect 5987 22276 5991 22332
rect 5927 22272 5991 22276
rect 6007 22332 6071 22336
rect 6007 22276 6011 22332
rect 6011 22276 6067 22332
rect 6067 22276 6071 22332
rect 6007 22272 6071 22276
rect 6087 22332 6151 22336
rect 6087 22276 6091 22332
rect 6091 22276 6147 22332
rect 6147 22276 6151 22332
rect 6087 22272 6151 22276
rect 9111 22332 9175 22336
rect 9111 22276 9115 22332
rect 9115 22276 9171 22332
rect 9171 22276 9175 22332
rect 9111 22272 9175 22276
rect 9191 22332 9255 22336
rect 9191 22276 9195 22332
rect 9195 22276 9251 22332
rect 9251 22276 9255 22332
rect 9191 22272 9255 22276
rect 9271 22332 9335 22336
rect 9271 22276 9275 22332
rect 9275 22276 9331 22332
rect 9331 22276 9335 22332
rect 9271 22272 9335 22276
rect 9351 22332 9415 22336
rect 9351 22276 9355 22332
rect 9355 22276 9411 22332
rect 9411 22276 9415 22332
rect 9351 22272 9415 22276
rect 4215 21788 4279 21792
rect 4215 21732 4219 21788
rect 4219 21732 4275 21788
rect 4275 21732 4279 21788
rect 4215 21728 4279 21732
rect 4295 21788 4359 21792
rect 4295 21732 4299 21788
rect 4299 21732 4355 21788
rect 4355 21732 4359 21788
rect 4295 21728 4359 21732
rect 4375 21788 4439 21792
rect 4375 21732 4379 21788
rect 4379 21732 4435 21788
rect 4435 21732 4439 21788
rect 4375 21728 4439 21732
rect 4455 21788 4519 21792
rect 4455 21732 4459 21788
rect 4459 21732 4515 21788
rect 4515 21732 4519 21788
rect 4455 21728 4519 21732
rect 7479 21788 7543 21792
rect 7479 21732 7483 21788
rect 7483 21732 7539 21788
rect 7539 21732 7543 21788
rect 7479 21728 7543 21732
rect 7559 21788 7623 21792
rect 7559 21732 7563 21788
rect 7563 21732 7619 21788
rect 7619 21732 7623 21788
rect 7559 21728 7623 21732
rect 7639 21788 7703 21792
rect 7639 21732 7643 21788
rect 7643 21732 7699 21788
rect 7699 21732 7703 21788
rect 7639 21728 7703 21732
rect 7719 21788 7783 21792
rect 7719 21732 7723 21788
rect 7723 21732 7779 21788
rect 7779 21732 7783 21788
rect 7719 21728 7783 21732
rect 2584 21244 2648 21248
rect 2584 21188 2588 21244
rect 2588 21188 2644 21244
rect 2644 21188 2648 21244
rect 2584 21184 2648 21188
rect 2664 21244 2728 21248
rect 2664 21188 2668 21244
rect 2668 21188 2724 21244
rect 2724 21188 2728 21244
rect 2664 21184 2728 21188
rect 2744 21244 2808 21248
rect 2744 21188 2748 21244
rect 2748 21188 2804 21244
rect 2804 21188 2808 21244
rect 2744 21184 2808 21188
rect 2824 21244 2888 21248
rect 2824 21188 2828 21244
rect 2828 21188 2884 21244
rect 2884 21188 2888 21244
rect 2824 21184 2888 21188
rect 5847 21244 5911 21248
rect 5847 21188 5851 21244
rect 5851 21188 5907 21244
rect 5907 21188 5911 21244
rect 5847 21184 5911 21188
rect 5927 21244 5991 21248
rect 5927 21188 5931 21244
rect 5931 21188 5987 21244
rect 5987 21188 5991 21244
rect 5927 21184 5991 21188
rect 6007 21244 6071 21248
rect 6007 21188 6011 21244
rect 6011 21188 6067 21244
rect 6067 21188 6071 21244
rect 6007 21184 6071 21188
rect 6087 21244 6151 21248
rect 6087 21188 6091 21244
rect 6091 21188 6147 21244
rect 6147 21188 6151 21244
rect 6087 21184 6151 21188
rect 9111 21244 9175 21248
rect 9111 21188 9115 21244
rect 9115 21188 9171 21244
rect 9171 21188 9175 21244
rect 9111 21184 9175 21188
rect 9191 21244 9255 21248
rect 9191 21188 9195 21244
rect 9195 21188 9251 21244
rect 9251 21188 9255 21244
rect 9191 21184 9255 21188
rect 9271 21244 9335 21248
rect 9271 21188 9275 21244
rect 9275 21188 9331 21244
rect 9331 21188 9335 21244
rect 9271 21184 9335 21188
rect 9351 21244 9415 21248
rect 9351 21188 9355 21244
rect 9355 21188 9411 21244
rect 9411 21188 9415 21244
rect 9351 21184 9415 21188
rect 4215 20700 4279 20704
rect 4215 20644 4219 20700
rect 4219 20644 4275 20700
rect 4275 20644 4279 20700
rect 4215 20640 4279 20644
rect 4295 20700 4359 20704
rect 4295 20644 4299 20700
rect 4299 20644 4355 20700
rect 4355 20644 4359 20700
rect 4295 20640 4359 20644
rect 4375 20700 4439 20704
rect 4375 20644 4379 20700
rect 4379 20644 4435 20700
rect 4435 20644 4439 20700
rect 4375 20640 4439 20644
rect 4455 20700 4519 20704
rect 4455 20644 4459 20700
rect 4459 20644 4515 20700
rect 4515 20644 4519 20700
rect 4455 20640 4519 20644
rect 7479 20700 7543 20704
rect 7479 20644 7483 20700
rect 7483 20644 7539 20700
rect 7539 20644 7543 20700
rect 7479 20640 7543 20644
rect 7559 20700 7623 20704
rect 7559 20644 7563 20700
rect 7563 20644 7619 20700
rect 7619 20644 7623 20700
rect 7559 20640 7623 20644
rect 7639 20700 7703 20704
rect 7639 20644 7643 20700
rect 7643 20644 7699 20700
rect 7699 20644 7703 20700
rect 7639 20640 7703 20644
rect 7719 20700 7783 20704
rect 7719 20644 7723 20700
rect 7723 20644 7779 20700
rect 7779 20644 7783 20700
rect 7719 20640 7783 20644
rect 2584 20156 2648 20160
rect 2584 20100 2588 20156
rect 2588 20100 2644 20156
rect 2644 20100 2648 20156
rect 2584 20096 2648 20100
rect 2664 20156 2728 20160
rect 2664 20100 2668 20156
rect 2668 20100 2724 20156
rect 2724 20100 2728 20156
rect 2664 20096 2728 20100
rect 2744 20156 2808 20160
rect 2744 20100 2748 20156
rect 2748 20100 2804 20156
rect 2804 20100 2808 20156
rect 2744 20096 2808 20100
rect 2824 20156 2888 20160
rect 2824 20100 2828 20156
rect 2828 20100 2884 20156
rect 2884 20100 2888 20156
rect 2824 20096 2888 20100
rect 5847 20156 5911 20160
rect 5847 20100 5851 20156
rect 5851 20100 5907 20156
rect 5907 20100 5911 20156
rect 5847 20096 5911 20100
rect 5927 20156 5991 20160
rect 5927 20100 5931 20156
rect 5931 20100 5987 20156
rect 5987 20100 5991 20156
rect 5927 20096 5991 20100
rect 6007 20156 6071 20160
rect 6007 20100 6011 20156
rect 6011 20100 6067 20156
rect 6067 20100 6071 20156
rect 6007 20096 6071 20100
rect 6087 20156 6151 20160
rect 6087 20100 6091 20156
rect 6091 20100 6147 20156
rect 6147 20100 6151 20156
rect 6087 20096 6151 20100
rect 9111 20156 9175 20160
rect 9111 20100 9115 20156
rect 9115 20100 9171 20156
rect 9171 20100 9175 20156
rect 9111 20096 9175 20100
rect 9191 20156 9255 20160
rect 9191 20100 9195 20156
rect 9195 20100 9251 20156
rect 9251 20100 9255 20156
rect 9191 20096 9255 20100
rect 9271 20156 9335 20160
rect 9271 20100 9275 20156
rect 9275 20100 9331 20156
rect 9331 20100 9335 20156
rect 9271 20096 9335 20100
rect 9351 20156 9415 20160
rect 9351 20100 9355 20156
rect 9355 20100 9411 20156
rect 9411 20100 9415 20156
rect 9351 20096 9415 20100
rect 4215 19612 4279 19616
rect 4215 19556 4219 19612
rect 4219 19556 4275 19612
rect 4275 19556 4279 19612
rect 4215 19552 4279 19556
rect 4295 19612 4359 19616
rect 4295 19556 4299 19612
rect 4299 19556 4355 19612
rect 4355 19556 4359 19612
rect 4295 19552 4359 19556
rect 4375 19612 4439 19616
rect 4375 19556 4379 19612
rect 4379 19556 4435 19612
rect 4435 19556 4439 19612
rect 4375 19552 4439 19556
rect 4455 19612 4519 19616
rect 4455 19556 4459 19612
rect 4459 19556 4515 19612
rect 4515 19556 4519 19612
rect 4455 19552 4519 19556
rect 7479 19612 7543 19616
rect 7479 19556 7483 19612
rect 7483 19556 7539 19612
rect 7539 19556 7543 19612
rect 7479 19552 7543 19556
rect 7559 19612 7623 19616
rect 7559 19556 7563 19612
rect 7563 19556 7619 19612
rect 7619 19556 7623 19612
rect 7559 19552 7623 19556
rect 7639 19612 7703 19616
rect 7639 19556 7643 19612
rect 7643 19556 7699 19612
rect 7699 19556 7703 19612
rect 7639 19552 7703 19556
rect 7719 19612 7783 19616
rect 7719 19556 7723 19612
rect 7723 19556 7779 19612
rect 7779 19556 7783 19612
rect 7719 19552 7783 19556
rect 2584 19068 2648 19072
rect 2584 19012 2588 19068
rect 2588 19012 2644 19068
rect 2644 19012 2648 19068
rect 2584 19008 2648 19012
rect 2664 19068 2728 19072
rect 2664 19012 2668 19068
rect 2668 19012 2724 19068
rect 2724 19012 2728 19068
rect 2664 19008 2728 19012
rect 2744 19068 2808 19072
rect 2744 19012 2748 19068
rect 2748 19012 2804 19068
rect 2804 19012 2808 19068
rect 2744 19008 2808 19012
rect 2824 19068 2888 19072
rect 2824 19012 2828 19068
rect 2828 19012 2884 19068
rect 2884 19012 2888 19068
rect 2824 19008 2888 19012
rect 5847 19068 5911 19072
rect 5847 19012 5851 19068
rect 5851 19012 5907 19068
rect 5907 19012 5911 19068
rect 5847 19008 5911 19012
rect 5927 19068 5991 19072
rect 5927 19012 5931 19068
rect 5931 19012 5987 19068
rect 5987 19012 5991 19068
rect 5927 19008 5991 19012
rect 6007 19068 6071 19072
rect 6007 19012 6011 19068
rect 6011 19012 6067 19068
rect 6067 19012 6071 19068
rect 6007 19008 6071 19012
rect 6087 19068 6151 19072
rect 6087 19012 6091 19068
rect 6091 19012 6147 19068
rect 6147 19012 6151 19068
rect 6087 19008 6151 19012
rect 9111 19068 9175 19072
rect 9111 19012 9115 19068
rect 9115 19012 9171 19068
rect 9171 19012 9175 19068
rect 9111 19008 9175 19012
rect 9191 19068 9255 19072
rect 9191 19012 9195 19068
rect 9195 19012 9251 19068
rect 9251 19012 9255 19068
rect 9191 19008 9255 19012
rect 9271 19068 9335 19072
rect 9271 19012 9275 19068
rect 9275 19012 9331 19068
rect 9331 19012 9335 19068
rect 9271 19008 9335 19012
rect 9351 19068 9415 19072
rect 9351 19012 9355 19068
rect 9355 19012 9411 19068
rect 9411 19012 9415 19068
rect 9351 19008 9415 19012
rect 4215 18524 4279 18528
rect 4215 18468 4219 18524
rect 4219 18468 4275 18524
rect 4275 18468 4279 18524
rect 4215 18464 4279 18468
rect 4295 18524 4359 18528
rect 4295 18468 4299 18524
rect 4299 18468 4355 18524
rect 4355 18468 4359 18524
rect 4295 18464 4359 18468
rect 4375 18524 4439 18528
rect 4375 18468 4379 18524
rect 4379 18468 4435 18524
rect 4435 18468 4439 18524
rect 4375 18464 4439 18468
rect 4455 18524 4519 18528
rect 4455 18468 4459 18524
rect 4459 18468 4515 18524
rect 4515 18468 4519 18524
rect 4455 18464 4519 18468
rect 7479 18524 7543 18528
rect 7479 18468 7483 18524
rect 7483 18468 7539 18524
rect 7539 18468 7543 18524
rect 7479 18464 7543 18468
rect 7559 18524 7623 18528
rect 7559 18468 7563 18524
rect 7563 18468 7619 18524
rect 7619 18468 7623 18524
rect 7559 18464 7623 18468
rect 7639 18524 7703 18528
rect 7639 18468 7643 18524
rect 7643 18468 7699 18524
rect 7699 18468 7703 18524
rect 7639 18464 7703 18468
rect 7719 18524 7783 18528
rect 7719 18468 7723 18524
rect 7723 18468 7779 18524
rect 7779 18468 7783 18524
rect 7719 18464 7783 18468
rect 2584 17980 2648 17984
rect 2584 17924 2588 17980
rect 2588 17924 2644 17980
rect 2644 17924 2648 17980
rect 2584 17920 2648 17924
rect 2664 17980 2728 17984
rect 2664 17924 2668 17980
rect 2668 17924 2724 17980
rect 2724 17924 2728 17980
rect 2664 17920 2728 17924
rect 2744 17980 2808 17984
rect 2744 17924 2748 17980
rect 2748 17924 2804 17980
rect 2804 17924 2808 17980
rect 2744 17920 2808 17924
rect 2824 17980 2888 17984
rect 2824 17924 2828 17980
rect 2828 17924 2884 17980
rect 2884 17924 2888 17980
rect 2824 17920 2888 17924
rect 5847 17980 5911 17984
rect 5847 17924 5851 17980
rect 5851 17924 5907 17980
rect 5907 17924 5911 17980
rect 5847 17920 5911 17924
rect 5927 17980 5991 17984
rect 5927 17924 5931 17980
rect 5931 17924 5987 17980
rect 5987 17924 5991 17980
rect 5927 17920 5991 17924
rect 6007 17980 6071 17984
rect 6007 17924 6011 17980
rect 6011 17924 6067 17980
rect 6067 17924 6071 17980
rect 6007 17920 6071 17924
rect 6087 17980 6151 17984
rect 6087 17924 6091 17980
rect 6091 17924 6147 17980
rect 6147 17924 6151 17980
rect 6087 17920 6151 17924
rect 9111 17980 9175 17984
rect 9111 17924 9115 17980
rect 9115 17924 9171 17980
rect 9171 17924 9175 17980
rect 9111 17920 9175 17924
rect 9191 17980 9255 17984
rect 9191 17924 9195 17980
rect 9195 17924 9251 17980
rect 9251 17924 9255 17980
rect 9191 17920 9255 17924
rect 9271 17980 9335 17984
rect 9271 17924 9275 17980
rect 9275 17924 9331 17980
rect 9331 17924 9335 17980
rect 9271 17920 9335 17924
rect 9351 17980 9415 17984
rect 9351 17924 9355 17980
rect 9355 17924 9411 17980
rect 9411 17924 9415 17980
rect 9351 17920 9415 17924
rect 4215 17436 4279 17440
rect 4215 17380 4219 17436
rect 4219 17380 4275 17436
rect 4275 17380 4279 17436
rect 4215 17376 4279 17380
rect 4295 17436 4359 17440
rect 4295 17380 4299 17436
rect 4299 17380 4355 17436
rect 4355 17380 4359 17436
rect 4295 17376 4359 17380
rect 4375 17436 4439 17440
rect 4375 17380 4379 17436
rect 4379 17380 4435 17436
rect 4435 17380 4439 17436
rect 4375 17376 4439 17380
rect 4455 17436 4519 17440
rect 4455 17380 4459 17436
rect 4459 17380 4515 17436
rect 4515 17380 4519 17436
rect 4455 17376 4519 17380
rect 7479 17436 7543 17440
rect 7479 17380 7483 17436
rect 7483 17380 7539 17436
rect 7539 17380 7543 17436
rect 7479 17376 7543 17380
rect 7559 17436 7623 17440
rect 7559 17380 7563 17436
rect 7563 17380 7619 17436
rect 7619 17380 7623 17436
rect 7559 17376 7623 17380
rect 7639 17436 7703 17440
rect 7639 17380 7643 17436
rect 7643 17380 7699 17436
rect 7699 17380 7703 17436
rect 7639 17376 7703 17380
rect 7719 17436 7783 17440
rect 7719 17380 7723 17436
rect 7723 17380 7779 17436
rect 7779 17380 7783 17436
rect 7719 17376 7783 17380
rect 2584 16892 2648 16896
rect 2584 16836 2588 16892
rect 2588 16836 2644 16892
rect 2644 16836 2648 16892
rect 2584 16832 2648 16836
rect 2664 16892 2728 16896
rect 2664 16836 2668 16892
rect 2668 16836 2724 16892
rect 2724 16836 2728 16892
rect 2664 16832 2728 16836
rect 2744 16892 2808 16896
rect 2744 16836 2748 16892
rect 2748 16836 2804 16892
rect 2804 16836 2808 16892
rect 2744 16832 2808 16836
rect 2824 16892 2888 16896
rect 2824 16836 2828 16892
rect 2828 16836 2884 16892
rect 2884 16836 2888 16892
rect 2824 16832 2888 16836
rect 5847 16892 5911 16896
rect 5847 16836 5851 16892
rect 5851 16836 5907 16892
rect 5907 16836 5911 16892
rect 5847 16832 5911 16836
rect 5927 16892 5991 16896
rect 5927 16836 5931 16892
rect 5931 16836 5987 16892
rect 5987 16836 5991 16892
rect 5927 16832 5991 16836
rect 6007 16892 6071 16896
rect 6007 16836 6011 16892
rect 6011 16836 6067 16892
rect 6067 16836 6071 16892
rect 6007 16832 6071 16836
rect 6087 16892 6151 16896
rect 6087 16836 6091 16892
rect 6091 16836 6147 16892
rect 6147 16836 6151 16892
rect 6087 16832 6151 16836
rect 9111 16892 9175 16896
rect 9111 16836 9115 16892
rect 9115 16836 9171 16892
rect 9171 16836 9175 16892
rect 9111 16832 9175 16836
rect 9191 16892 9255 16896
rect 9191 16836 9195 16892
rect 9195 16836 9251 16892
rect 9251 16836 9255 16892
rect 9191 16832 9255 16836
rect 9271 16892 9335 16896
rect 9271 16836 9275 16892
rect 9275 16836 9331 16892
rect 9331 16836 9335 16892
rect 9271 16832 9335 16836
rect 9351 16892 9415 16896
rect 9351 16836 9355 16892
rect 9355 16836 9411 16892
rect 9411 16836 9415 16892
rect 9351 16832 9415 16836
rect 4215 16348 4279 16352
rect 4215 16292 4219 16348
rect 4219 16292 4275 16348
rect 4275 16292 4279 16348
rect 4215 16288 4279 16292
rect 4295 16348 4359 16352
rect 4295 16292 4299 16348
rect 4299 16292 4355 16348
rect 4355 16292 4359 16348
rect 4295 16288 4359 16292
rect 4375 16348 4439 16352
rect 4375 16292 4379 16348
rect 4379 16292 4435 16348
rect 4435 16292 4439 16348
rect 4375 16288 4439 16292
rect 4455 16348 4519 16352
rect 4455 16292 4459 16348
rect 4459 16292 4515 16348
rect 4515 16292 4519 16348
rect 4455 16288 4519 16292
rect 7479 16348 7543 16352
rect 7479 16292 7483 16348
rect 7483 16292 7539 16348
rect 7539 16292 7543 16348
rect 7479 16288 7543 16292
rect 7559 16348 7623 16352
rect 7559 16292 7563 16348
rect 7563 16292 7619 16348
rect 7619 16292 7623 16348
rect 7559 16288 7623 16292
rect 7639 16348 7703 16352
rect 7639 16292 7643 16348
rect 7643 16292 7699 16348
rect 7699 16292 7703 16348
rect 7639 16288 7703 16292
rect 7719 16348 7783 16352
rect 7719 16292 7723 16348
rect 7723 16292 7779 16348
rect 7779 16292 7783 16348
rect 7719 16288 7783 16292
rect 2584 15804 2648 15808
rect 2584 15748 2588 15804
rect 2588 15748 2644 15804
rect 2644 15748 2648 15804
rect 2584 15744 2648 15748
rect 2664 15804 2728 15808
rect 2664 15748 2668 15804
rect 2668 15748 2724 15804
rect 2724 15748 2728 15804
rect 2664 15744 2728 15748
rect 2744 15804 2808 15808
rect 2744 15748 2748 15804
rect 2748 15748 2804 15804
rect 2804 15748 2808 15804
rect 2744 15744 2808 15748
rect 2824 15804 2888 15808
rect 2824 15748 2828 15804
rect 2828 15748 2884 15804
rect 2884 15748 2888 15804
rect 2824 15744 2888 15748
rect 5847 15804 5911 15808
rect 5847 15748 5851 15804
rect 5851 15748 5907 15804
rect 5907 15748 5911 15804
rect 5847 15744 5911 15748
rect 5927 15804 5991 15808
rect 5927 15748 5931 15804
rect 5931 15748 5987 15804
rect 5987 15748 5991 15804
rect 5927 15744 5991 15748
rect 6007 15804 6071 15808
rect 6007 15748 6011 15804
rect 6011 15748 6067 15804
rect 6067 15748 6071 15804
rect 6007 15744 6071 15748
rect 6087 15804 6151 15808
rect 6087 15748 6091 15804
rect 6091 15748 6147 15804
rect 6147 15748 6151 15804
rect 6087 15744 6151 15748
rect 9111 15804 9175 15808
rect 9111 15748 9115 15804
rect 9115 15748 9171 15804
rect 9171 15748 9175 15804
rect 9111 15744 9175 15748
rect 9191 15804 9255 15808
rect 9191 15748 9195 15804
rect 9195 15748 9251 15804
rect 9251 15748 9255 15804
rect 9191 15744 9255 15748
rect 9271 15804 9335 15808
rect 9271 15748 9275 15804
rect 9275 15748 9331 15804
rect 9331 15748 9335 15804
rect 9271 15744 9335 15748
rect 9351 15804 9415 15808
rect 9351 15748 9355 15804
rect 9355 15748 9411 15804
rect 9411 15748 9415 15804
rect 9351 15744 9415 15748
rect 4215 15260 4279 15264
rect 4215 15204 4219 15260
rect 4219 15204 4275 15260
rect 4275 15204 4279 15260
rect 4215 15200 4279 15204
rect 4295 15260 4359 15264
rect 4295 15204 4299 15260
rect 4299 15204 4355 15260
rect 4355 15204 4359 15260
rect 4295 15200 4359 15204
rect 4375 15260 4439 15264
rect 4375 15204 4379 15260
rect 4379 15204 4435 15260
rect 4435 15204 4439 15260
rect 4375 15200 4439 15204
rect 4455 15260 4519 15264
rect 4455 15204 4459 15260
rect 4459 15204 4515 15260
rect 4515 15204 4519 15260
rect 4455 15200 4519 15204
rect 7479 15260 7543 15264
rect 7479 15204 7483 15260
rect 7483 15204 7539 15260
rect 7539 15204 7543 15260
rect 7479 15200 7543 15204
rect 7559 15260 7623 15264
rect 7559 15204 7563 15260
rect 7563 15204 7619 15260
rect 7619 15204 7623 15260
rect 7559 15200 7623 15204
rect 7639 15260 7703 15264
rect 7639 15204 7643 15260
rect 7643 15204 7699 15260
rect 7699 15204 7703 15260
rect 7639 15200 7703 15204
rect 7719 15260 7783 15264
rect 7719 15204 7723 15260
rect 7723 15204 7779 15260
rect 7779 15204 7783 15260
rect 7719 15200 7783 15204
rect 2584 14716 2648 14720
rect 2584 14660 2588 14716
rect 2588 14660 2644 14716
rect 2644 14660 2648 14716
rect 2584 14656 2648 14660
rect 2664 14716 2728 14720
rect 2664 14660 2668 14716
rect 2668 14660 2724 14716
rect 2724 14660 2728 14716
rect 2664 14656 2728 14660
rect 2744 14716 2808 14720
rect 2744 14660 2748 14716
rect 2748 14660 2804 14716
rect 2804 14660 2808 14716
rect 2744 14656 2808 14660
rect 2824 14716 2888 14720
rect 2824 14660 2828 14716
rect 2828 14660 2884 14716
rect 2884 14660 2888 14716
rect 2824 14656 2888 14660
rect 5847 14716 5911 14720
rect 5847 14660 5851 14716
rect 5851 14660 5907 14716
rect 5907 14660 5911 14716
rect 5847 14656 5911 14660
rect 5927 14716 5991 14720
rect 5927 14660 5931 14716
rect 5931 14660 5987 14716
rect 5987 14660 5991 14716
rect 5927 14656 5991 14660
rect 6007 14716 6071 14720
rect 6007 14660 6011 14716
rect 6011 14660 6067 14716
rect 6067 14660 6071 14716
rect 6007 14656 6071 14660
rect 6087 14716 6151 14720
rect 6087 14660 6091 14716
rect 6091 14660 6147 14716
rect 6147 14660 6151 14716
rect 6087 14656 6151 14660
rect 9111 14716 9175 14720
rect 9111 14660 9115 14716
rect 9115 14660 9171 14716
rect 9171 14660 9175 14716
rect 9111 14656 9175 14660
rect 9191 14716 9255 14720
rect 9191 14660 9195 14716
rect 9195 14660 9251 14716
rect 9251 14660 9255 14716
rect 9191 14656 9255 14660
rect 9271 14716 9335 14720
rect 9271 14660 9275 14716
rect 9275 14660 9331 14716
rect 9331 14660 9335 14716
rect 9271 14656 9335 14660
rect 9351 14716 9415 14720
rect 9351 14660 9355 14716
rect 9355 14660 9411 14716
rect 9411 14660 9415 14716
rect 9351 14656 9415 14660
rect 4215 14172 4279 14176
rect 4215 14116 4219 14172
rect 4219 14116 4275 14172
rect 4275 14116 4279 14172
rect 4215 14112 4279 14116
rect 4295 14172 4359 14176
rect 4295 14116 4299 14172
rect 4299 14116 4355 14172
rect 4355 14116 4359 14172
rect 4295 14112 4359 14116
rect 4375 14172 4439 14176
rect 4375 14116 4379 14172
rect 4379 14116 4435 14172
rect 4435 14116 4439 14172
rect 4375 14112 4439 14116
rect 4455 14172 4519 14176
rect 4455 14116 4459 14172
rect 4459 14116 4515 14172
rect 4515 14116 4519 14172
rect 4455 14112 4519 14116
rect 7479 14172 7543 14176
rect 7479 14116 7483 14172
rect 7483 14116 7539 14172
rect 7539 14116 7543 14172
rect 7479 14112 7543 14116
rect 7559 14172 7623 14176
rect 7559 14116 7563 14172
rect 7563 14116 7619 14172
rect 7619 14116 7623 14172
rect 7559 14112 7623 14116
rect 7639 14172 7703 14176
rect 7639 14116 7643 14172
rect 7643 14116 7699 14172
rect 7699 14116 7703 14172
rect 7639 14112 7703 14116
rect 7719 14172 7783 14176
rect 7719 14116 7723 14172
rect 7723 14116 7779 14172
rect 7779 14116 7783 14172
rect 7719 14112 7783 14116
rect 2584 13628 2648 13632
rect 2584 13572 2588 13628
rect 2588 13572 2644 13628
rect 2644 13572 2648 13628
rect 2584 13568 2648 13572
rect 2664 13628 2728 13632
rect 2664 13572 2668 13628
rect 2668 13572 2724 13628
rect 2724 13572 2728 13628
rect 2664 13568 2728 13572
rect 2744 13628 2808 13632
rect 2744 13572 2748 13628
rect 2748 13572 2804 13628
rect 2804 13572 2808 13628
rect 2744 13568 2808 13572
rect 2824 13628 2888 13632
rect 2824 13572 2828 13628
rect 2828 13572 2884 13628
rect 2884 13572 2888 13628
rect 2824 13568 2888 13572
rect 5847 13628 5911 13632
rect 5847 13572 5851 13628
rect 5851 13572 5907 13628
rect 5907 13572 5911 13628
rect 5847 13568 5911 13572
rect 5927 13628 5991 13632
rect 5927 13572 5931 13628
rect 5931 13572 5987 13628
rect 5987 13572 5991 13628
rect 5927 13568 5991 13572
rect 6007 13628 6071 13632
rect 6007 13572 6011 13628
rect 6011 13572 6067 13628
rect 6067 13572 6071 13628
rect 6007 13568 6071 13572
rect 6087 13628 6151 13632
rect 6087 13572 6091 13628
rect 6091 13572 6147 13628
rect 6147 13572 6151 13628
rect 6087 13568 6151 13572
rect 9111 13628 9175 13632
rect 9111 13572 9115 13628
rect 9115 13572 9171 13628
rect 9171 13572 9175 13628
rect 9111 13568 9175 13572
rect 9191 13628 9255 13632
rect 9191 13572 9195 13628
rect 9195 13572 9251 13628
rect 9251 13572 9255 13628
rect 9191 13568 9255 13572
rect 9271 13628 9335 13632
rect 9271 13572 9275 13628
rect 9275 13572 9331 13628
rect 9331 13572 9335 13628
rect 9271 13568 9335 13572
rect 9351 13628 9415 13632
rect 9351 13572 9355 13628
rect 9355 13572 9411 13628
rect 9411 13572 9415 13628
rect 9351 13568 9415 13572
rect 4215 13084 4279 13088
rect 4215 13028 4219 13084
rect 4219 13028 4275 13084
rect 4275 13028 4279 13084
rect 4215 13024 4279 13028
rect 4295 13084 4359 13088
rect 4295 13028 4299 13084
rect 4299 13028 4355 13084
rect 4355 13028 4359 13084
rect 4295 13024 4359 13028
rect 4375 13084 4439 13088
rect 4375 13028 4379 13084
rect 4379 13028 4435 13084
rect 4435 13028 4439 13084
rect 4375 13024 4439 13028
rect 4455 13084 4519 13088
rect 4455 13028 4459 13084
rect 4459 13028 4515 13084
rect 4515 13028 4519 13084
rect 4455 13024 4519 13028
rect 7479 13084 7543 13088
rect 7479 13028 7483 13084
rect 7483 13028 7539 13084
rect 7539 13028 7543 13084
rect 7479 13024 7543 13028
rect 7559 13084 7623 13088
rect 7559 13028 7563 13084
rect 7563 13028 7619 13084
rect 7619 13028 7623 13084
rect 7559 13024 7623 13028
rect 7639 13084 7703 13088
rect 7639 13028 7643 13084
rect 7643 13028 7699 13084
rect 7699 13028 7703 13084
rect 7639 13024 7703 13028
rect 7719 13084 7783 13088
rect 7719 13028 7723 13084
rect 7723 13028 7779 13084
rect 7779 13028 7783 13084
rect 7719 13024 7783 13028
rect 2584 12540 2648 12544
rect 2584 12484 2588 12540
rect 2588 12484 2644 12540
rect 2644 12484 2648 12540
rect 2584 12480 2648 12484
rect 2664 12540 2728 12544
rect 2664 12484 2668 12540
rect 2668 12484 2724 12540
rect 2724 12484 2728 12540
rect 2664 12480 2728 12484
rect 2744 12540 2808 12544
rect 2744 12484 2748 12540
rect 2748 12484 2804 12540
rect 2804 12484 2808 12540
rect 2744 12480 2808 12484
rect 2824 12540 2888 12544
rect 2824 12484 2828 12540
rect 2828 12484 2884 12540
rect 2884 12484 2888 12540
rect 2824 12480 2888 12484
rect 5847 12540 5911 12544
rect 5847 12484 5851 12540
rect 5851 12484 5907 12540
rect 5907 12484 5911 12540
rect 5847 12480 5911 12484
rect 5927 12540 5991 12544
rect 5927 12484 5931 12540
rect 5931 12484 5987 12540
rect 5987 12484 5991 12540
rect 5927 12480 5991 12484
rect 6007 12540 6071 12544
rect 6007 12484 6011 12540
rect 6011 12484 6067 12540
rect 6067 12484 6071 12540
rect 6007 12480 6071 12484
rect 6087 12540 6151 12544
rect 6087 12484 6091 12540
rect 6091 12484 6147 12540
rect 6147 12484 6151 12540
rect 6087 12480 6151 12484
rect 9111 12540 9175 12544
rect 9111 12484 9115 12540
rect 9115 12484 9171 12540
rect 9171 12484 9175 12540
rect 9111 12480 9175 12484
rect 9191 12540 9255 12544
rect 9191 12484 9195 12540
rect 9195 12484 9251 12540
rect 9251 12484 9255 12540
rect 9191 12480 9255 12484
rect 9271 12540 9335 12544
rect 9271 12484 9275 12540
rect 9275 12484 9331 12540
rect 9331 12484 9335 12540
rect 9271 12480 9335 12484
rect 9351 12540 9415 12544
rect 9351 12484 9355 12540
rect 9355 12484 9411 12540
rect 9411 12484 9415 12540
rect 9351 12480 9415 12484
rect 4215 11996 4279 12000
rect 4215 11940 4219 11996
rect 4219 11940 4275 11996
rect 4275 11940 4279 11996
rect 4215 11936 4279 11940
rect 4295 11996 4359 12000
rect 4295 11940 4299 11996
rect 4299 11940 4355 11996
rect 4355 11940 4359 11996
rect 4295 11936 4359 11940
rect 4375 11996 4439 12000
rect 4375 11940 4379 11996
rect 4379 11940 4435 11996
rect 4435 11940 4439 11996
rect 4375 11936 4439 11940
rect 4455 11996 4519 12000
rect 4455 11940 4459 11996
rect 4459 11940 4515 11996
rect 4515 11940 4519 11996
rect 4455 11936 4519 11940
rect 7479 11996 7543 12000
rect 7479 11940 7483 11996
rect 7483 11940 7539 11996
rect 7539 11940 7543 11996
rect 7479 11936 7543 11940
rect 7559 11996 7623 12000
rect 7559 11940 7563 11996
rect 7563 11940 7619 11996
rect 7619 11940 7623 11996
rect 7559 11936 7623 11940
rect 7639 11996 7703 12000
rect 7639 11940 7643 11996
rect 7643 11940 7699 11996
rect 7699 11940 7703 11996
rect 7639 11936 7703 11940
rect 7719 11996 7783 12000
rect 7719 11940 7723 11996
rect 7723 11940 7779 11996
rect 7779 11940 7783 11996
rect 7719 11936 7783 11940
rect 2584 11452 2648 11456
rect 2584 11396 2588 11452
rect 2588 11396 2644 11452
rect 2644 11396 2648 11452
rect 2584 11392 2648 11396
rect 2664 11452 2728 11456
rect 2664 11396 2668 11452
rect 2668 11396 2724 11452
rect 2724 11396 2728 11452
rect 2664 11392 2728 11396
rect 2744 11452 2808 11456
rect 2744 11396 2748 11452
rect 2748 11396 2804 11452
rect 2804 11396 2808 11452
rect 2744 11392 2808 11396
rect 2824 11452 2888 11456
rect 2824 11396 2828 11452
rect 2828 11396 2884 11452
rect 2884 11396 2888 11452
rect 2824 11392 2888 11396
rect 5847 11452 5911 11456
rect 5847 11396 5851 11452
rect 5851 11396 5907 11452
rect 5907 11396 5911 11452
rect 5847 11392 5911 11396
rect 5927 11452 5991 11456
rect 5927 11396 5931 11452
rect 5931 11396 5987 11452
rect 5987 11396 5991 11452
rect 5927 11392 5991 11396
rect 6007 11452 6071 11456
rect 6007 11396 6011 11452
rect 6011 11396 6067 11452
rect 6067 11396 6071 11452
rect 6007 11392 6071 11396
rect 6087 11452 6151 11456
rect 6087 11396 6091 11452
rect 6091 11396 6147 11452
rect 6147 11396 6151 11452
rect 6087 11392 6151 11396
rect 9111 11452 9175 11456
rect 9111 11396 9115 11452
rect 9115 11396 9171 11452
rect 9171 11396 9175 11452
rect 9111 11392 9175 11396
rect 9191 11452 9255 11456
rect 9191 11396 9195 11452
rect 9195 11396 9251 11452
rect 9251 11396 9255 11452
rect 9191 11392 9255 11396
rect 9271 11452 9335 11456
rect 9271 11396 9275 11452
rect 9275 11396 9331 11452
rect 9331 11396 9335 11452
rect 9271 11392 9335 11396
rect 9351 11452 9415 11456
rect 9351 11396 9355 11452
rect 9355 11396 9411 11452
rect 9411 11396 9415 11452
rect 9351 11392 9415 11396
rect 4215 10908 4279 10912
rect 4215 10852 4219 10908
rect 4219 10852 4275 10908
rect 4275 10852 4279 10908
rect 4215 10848 4279 10852
rect 4295 10908 4359 10912
rect 4295 10852 4299 10908
rect 4299 10852 4355 10908
rect 4355 10852 4359 10908
rect 4295 10848 4359 10852
rect 4375 10908 4439 10912
rect 4375 10852 4379 10908
rect 4379 10852 4435 10908
rect 4435 10852 4439 10908
rect 4375 10848 4439 10852
rect 4455 10908 4519 10912
rect 4455 10852 4459 10908
rect 4459 10852 4515 10908
rect 4515 10852 4519 10908
rect 4455 10848 4519 10852
rect 7479 10908 7543 10912
rect 7479 10852 7483 10908
rect 7483 10852 7539 10908
rect 7539 10852 7543 10908
rect 7479 10848 7543 10852
rect 7559 10908 7623 10912
rect 7559 10852 7563 10908
rect 7563 10852 7619 10908
rect 7619 10852 7623 10908
rect 7559 10848 7623 10852
rect 7639 10908 7703 10912
rect 7639 10852 7643 10908
rect 7643 10852 7699 10908
rect 7699 10852 7703 10908
rect 7639 10848 7703 10852
rect 7719 10908 7783 10912
rect 7719 10852 7723 10908
rect 7723 10852 7779 10908
rect 7779 10852 7783 10908
rect 7719 10848 7783 10852
rect 2584 10364 2648 10368
rect 2584 10308 2588 10364
rect 2588 10308 2644 10364
rect 2644 10308 2648 10364
rect 2584 10304 2648 10308
rect 2664 10364 2728 10368
rect 2664 10308 2668 10364
rect 2668 10308 2724 10364
rect 2724 10308 2728 10364
rect 2664 10304 2728 10308
rect 2744 10364 2808 10368
rect 2744 10308 2748 10364
rect 2748 10308 2804 10364
rect 2804 10308 2808 10364
rect 2744 10304 2808 10308
rect 2824 10364 2888 10368
rect 2824 10308 2828 10364
rect 2828 10308 2884 10364
rect 2884 10308 2888 10364
rect 2824 10304 2888 10308
rect 5847 10364 5911 10368
rect 5847 10308 5851 10364
rect 5851 10308 5907 10364
rect 5907 10308 5911 10364
rect 5847 10304 5911 10308
rect 5927 10364 5991 10368
rect 5927 10308 5931 10364
rect 5931 10308 5987 10364
rect 5987 10308 5991 10364
rect 5927 10304 5991 10308
rect 6007 10364 6071 10368
rect 6007 10308 6011 10364
rect 6011 10308 6067 10364
rect 6067 10308 6071 10364
rect 6007 10304 6071 10308
rect 6087 10364 6151 10368
rect 6087 10308 6091 10364
rect 6091 10308 6147 10364
rect 6147 10308 6151 10364
rect 6087 10304 6151 10308
rect 9111 10364 9175 10368
rect 9111 10308 9115 10364
rect 9115 10308 9171 10364
rect 9171 10308 9175 10364
rect 9111 10304 9175 10308
rect 9191 10364 9255 10368
rect 9191 10308 9195 10364
rect 9195 10308 9251 10364
rect 9251 10308 9255 10364
rect 9191 10304 9255 10308
rect 9271 10364 9335 10368
rect 9271 10308 9275 10364
rect 9275 10308 9331 10364
rect 9331 10308 9335 10364
rect 9271 10304 9335 10308
rect 9351 10364 9415 10368
rect 9351 10308 9355 10364
rect 9355 10308 9411 10364
rect 9411 10308 9415 10364
rect 9351 10304 9415 10308
rect 4215 9820 4279 9824
rect 4215 9764 4219 9820
rect 4219 9764 4275 9820
rect 4275 9764 4279 9820
rect 4215 9760 4279 9764
rect 4295 9820 4359 9824
rect 4295 9764 4299 9820
rect 4299 9764 4355 9820
rect 4355 9764 4359 9820
rect 4295 9760 4359 9764
rect 4375 9820 4439 9824
rect 4375 9764 4379 9820
rect 4379 9764 4435 9820
rect 4435 9764 4439 9820
rect 4375 9760 4439 9764
rect 4455 9820 4519 9824
rect 4455 9764 4459 9820
rect 4459 9764 4515 9820
rect 4515 9764 4519 9820
rect 4455 9760 4519 9764
rect 7479 9820 7543 9824
rect 7479 9764 7483 9820
rect 7483 9764 7539 9820
rect 7539 9764 7543 9820
rect 7479 9760 7543 9764
rect 7559 9820 7623 9824
rect 7559 9764 7563 9820
rect 7563 9764 7619 9820
rect 7619 9764 7623 9820
rect 7559 9760 7623 9764
rect 7639 9820 7703 9824
rect 7639 9764 7643 9820
rect 7643 9764 7699 9820
rect 7699 9764 7703 9820
rect 7639 9760 7703 9764
rect 7719 9820 7783 9824
rect 7719 9764 7723 9820
rect 7723 9764 7779 9820
rect 7779 9764 7783 9820
rect 7719 9760 7783 9764
rect 2584 9276 2648 9280
rect 2584 9220 2588 9276
rect 2588 9220 2644 9276
rect 2644 9220 2648 9276
rect 2584 9216 2648 9220
rect 2664 9276 2728 9280
rect 2664 9220 2668 9276
rect 2668 9220 2724 9276
rect 2724 9220 2728 9276
rect 2664 9216 2728 9220
rect 2744 9276 2808 9280
rect 2744 9220 2748 9276
rect 2748 9220 2804 9276
rect 2804 9220 2808 9276
rect 2744 9216 2808 9220
rect 2824 9276 2888 9280
rect 2824 9220 2828 9276
rect 2828 9220 2884 9276
rect 2884 9220 2888 9276
rect 2824 9216 2888 9220
rect 5847 9276 5911 9280
rect 5847 9220 5851 9276
rect 5851 9220 5907 9276
rect 5907 9220 5911 9276
rect 5847 9216 5911 9220
rect 5927 9276 5991 9280
rect 5927 9220 5931 9276
rect 5931 9220 5987 9276
rect 5987 9220 5991 9276
rect 5927 9216 5991 9220
rect 6007 9276 6071 9280
rect 6007 9220 6011 9276
rect 6011 9220 6067 9276
rect 6067 9220 6071 9276
rect 6007 9216 6071 9220
rect 6087 9276 6151 9280
rect 6087 9220 6091 9276
rect 6091 9220 6147 9276
rect 6147 9220 6151 9276
rect 6087 9216 6151 9220
rect 9111 9276 9175 9280
rect 9111 9220 9115 9276
rect 9115 9220 9171 9276
rect 9171 9220 9175 9276
rect 9111 9216 9175 9220
rect 9191 9276 9255 9280
rect 9191 9220 9195 9276
rect 9195 9220 9251 9276
rect 9251 9220 9255 9276
rect 9191 9216 9255 9220
rect 9271 9276 9335 9280
rect 9271 9220 9275 9276
rect 9275 9220 9331 9276
rect 9331 9220 9335 9276
rect 9271 9216 9335 9220
rect 9351 9276 9415 9280
rect 9351 9220 9355 9276
rect 9355 9220 9411 9276
rect 9411 9220 9415 9276
rect 9351 9216 9415 9220
rect 4215 8732 4279 8736
rect 4215 8676 4219 8732
rect 4219 8676 4275 8732
rect 4275 8676 4279 8732
rect 4215 8672 4279 8676
rect 4295 8732 4359 8736
rect 4295 8676 4299 8732
rect 4299 8676 4355 8732
rect 4355 8676 4359 8732
rect 4295 8672 4359 8676
rect 4375 8732 4439 8736
rect 4375 8676 4379 8732
rect 4379 8676 4435 8732
rect 4435 8676 4439 8732
rect 4375 8672 4439 8676
rect 4455 8732 4519 8736
rect 4455 8676 4459 8732
rect 4459 8676 4515 8732
rect 4515 8676 4519 8732
rect 4455 8672 4519 8676
rect 7479 8732 7543 8736
rect 7479 8676 7483 8732
rect 7483 8676 7539 8732
rect 7539 8676 7543 8732
rect 7479 8672 7543 8676
rect 7559 8732 7623 8736
rect 7559 8676 7563 8732
rect 7563 8676 7619 8732
rect 7619 8676 7623 8732
rect 7559 8672 7623 8676
rect 7639 8732 7703 8736
rect 7639 8676 7643 8732
rect 7643 8676 7699 8732
rect 7699 8676 7703 8732
rect 7639 8672 7703 8676
rect 7719 8732 7783 8736
rect 7719 8676 7723 8732
rect 7723 8676 7779 8732
rect 7779 8676 7783 8732
rect 7719 8672 7783 8676
rect 2584 8188 2648 8192
rect 2584 8132 2588 8188
rect 2588 8132 2644 8188
rect 2644 8132 2648 8188
rect 2584 8128 2648 8132
rect 2664 8188 2728 8192
rect 2664 8132 2668 8188
rect 2668 8132 2724 8188
rect 2724 8132 2728 8188
rect 2664 8128 2728 8132
rect 2744 8188 2808 8192
rect 2744 8132 2748 8188
rect 2748 8132 2804 8188
rect 2804 8132 2808 8188
rect 2744 8128 2808 8132
rect 2824 8188 2888 8192
rect 2824 8132 2828 8188
rect 2828 8132 2884 8188
rect 2884 8132 2888 8188
rect 2824 8128 2888 8132
rect 5847 8188 5911 8192
rect 5847 8132 5851 8188
rect 5851 8132 5907 8188
rect 5907 8132 5911 8188
rect 5847 8128 5911 8132
rect 5927 8188 5991 8192
rect 5927 8132 5931 8188
rect 5931 8132 5987 8188
rect 5987 8132 5991 8188
rect 5927 8128 5991 8132
rect 6007 8188 6071 8192
rect 6007 8132 6011 8188
rect 6011 8132 6067 8188
rect 6067 8132 6071 8188
rect 6007 8128 6071 8132
rect 6087 8188 6151 8192
rect 6087 8132 6091 8188
rect 6091 8132 6147 8188
rect 6147 8132 6151 8188
rect 6087 8128 6151 8132
rect 9111 8188 9175 8192
rect 9111 8132 9115 8188
rect 9115 8132 9171 8188
rect 9171 8132 9175 8188
rect 9111 8128 9175 8132
rect 9191 8188 9255 8192
rect 9191 8132 9195 8188
rect 9195 8132 9251 8188
rect 9251 8132 9255 8188
rect 9191 8128 9255 8132
rect 9271 8188 9335 8192
rect 9271 8132 9275 8188
rect 9275 8132 9331 8188
rect 9331 8132 9335 8188
rect 9271 8128 9335 8132
rect 9351 8188 9415 8192
rect 9351 8132 9355 8188
rect 9355 8132 9411 8188
rect 9411 8132 9415 8188
rect 9351 8128 9415 8132
rect 4215 7644 4279 7648
rect 4215 7588 4219 7644
rect 4219 7588 4275 7644
rect 4275 7588 4279 7644
rect 4215 7584 4279 7588
rect 4295 7644 4359 7648
rect 4295 7588 4299 7644
rect 4299 7588 4355 7644
rect 4355 7588 4359 7644
rect 4295 7584 4359 7588
rect 4375 7644 4439 7648
rect 4375 7588 4379 7644
rect 4379 7588 4435 7644
rect 4435 7588 4439 7644
rect 4375 7584 4439 7588
rect 4455 7644 4519 7648
rect 4455 7588 4459 7644
rect 4459 7588 4515 7644
rect 4515 7588 4519 7644
rect 4455 7584 4519 7588
rect 7479 7644 7543 7648
rect 7479 7588 7483 7644
rect 7483 7588 7539 7644
rect 7539 7588 7543 7644
rect 7479 7584 7543 7588
rect 7559 7644 7623 7648
rect 7559 7588 7563 7644
rect 7563 7588 7619 7644
rect 7619 7588 7623 7644
rect 7559 7584 7623 7588
rect 7639 7644 7703 7648
rect 7639 7588 7643 7644
rect 7643 7588 7699 7644
rect 7699 7588 7703 7644
rect 7639 7584 7703 7588
rect 7719 7644 7783 7648
rect 7719 7588 7723 7644
rect 7723 7588 7779 7644
rect 7779 7588 7783 7644
rect 7719 7584 7783 7588
rect 2584 7100 2648 7104
rect 2584 7044 2588 7100
rect 2588 7044 2644 7100
rect 2644 7044 2648 7100
rect 2584 7040 2648 7044
rect 2664 7100 2728 7104
rect 2664 7044 2668 7100
rect 2668 7044 2724 7100
rect 2724 7044 2728 7100
rect 2664 7040 2728 7044
rect 2744 7100 2808 7104
rect 2744 7044 2748 7100
rect 2748 7044 2804 7100
rect 2804 7044 2808 7100
rect 2744 7040 2808 7044
rect 2824 7100 2888 7104
rect 2824 7044 2828 7100
rect 2828 7044 2884 7100
rect 2884 7044 2888 7100
rect 2824 7040 2888 7044
rect 5847 7100 5911 7104
rect 5847 7044 5851 7100
rect 5851 7044 5907 7100
rect 5907 7044 5911 7100
rect 5847 7040 5911 7044
rect 5927 7100 5991 7104
rect 5927 7044 5931 7100
rect 5931 7044 5987 7100
rect 5987 7044 5991 7100
rect 5927 7040 5991 7044
rect 6007 7100 6071 7104
rect 6007 7044 6011 7100
rect 6011 7044 6067 7100
rect 6067 7044 6071 7100
rect 6007 7040 6071 7044
rect 6087 7100 6151 7104
rect 6087 7044 6091 7100
rect 6091 7044 6147 7100
rect 6147 7044 6151 7100
rect 6087 7040 6151 7044
rect 9111 7100 9175 7104
rect 9111 7044 9115 7100
rect 9115 7044 9171 7100
rect 9171 7044 9175 7100
rect 9111 7040 9175 7044
rect 9191 7100 9255 7104
rect 9191 7044 9195 7100
rect 9195 7044 9251 7100
rect 9251 7044 9255 7100
rect 9191 7040 9255 7044
rect 9271 7100 9335 7104
rect 9271 7044 9275 7100
rect 9275 7044 9331 7100
rect 9331 7044 9335 7100
rect 9271 7040 9335 7044
rect 9351 7100 9415 7104
rect 9351 7044 9355 7100
rect 9355 7044 9411 7100
rect 9411 7044 9415 7100
rect 9351 7040 9415 7044
rect 4215 6556 4279 6560
rect 4215 6500 4219 6556
rect 4219 6500 4275 6556
rect 4275 6500 4279 6556
rect 4215 6496 4279 6500
rect 4295 6556 4359 6560
rect 4295 6500 4299 6556
rect 4299 6500 4355 6556
rect 4355 6500 4359 6556
rect 4295 6496 4359 6500
rect 4375 6556 4439 6560
rect 4375 6500 4379 6556
rect 4379 6500 4435 6556
rect 4435 6500 4439 6556
rect 4375 6496 4439 6500
rect 4455 6556 4519 6560
rect 4455 6500 4459 6556
rect 4459 6500 4515 6556
rect 4515 6500 4519 6556
rect 4455 6496 4519 6500
rect 7479 6556 7543 6560
rect 7479 6500 7483 6556
rect 7483 6500 7539 6556
rect 7539 6500 7543 6556
rect 7479 6496 7543 6500
rect 7559 6556 7623 6560
rect 7559 6500 7563 6556
rect 7563 6500 7619 6556
rect 7619 6500 7623 6556
rect 7559 6496 7623 6500
rect 7639 6556 7703 6560
rect 7639 6500 7643 6556
rect 7643 6500 7699 6556
rect 7699 6500 7703 6556
rect 7639 6496 7703 6500
rect 7719 6556 7783 6560
rect 7719 6500 7723 6556
rect 7723 6500 7779 6556
rect 7779 6500 7783 6556
rect 7719 6496 7783 6500
rect 2584 6012 2648 6016
rect 2584 5956 2588 6012
rect 2588 5956 2644 6012
rect 2644 5956 2648 6012
rect 2584 5952 2648 5956
rect 2664 6012 2728 6016
rect 2664 5956 2668 6012
rect 2668 5956 2724 6012
rect 2724 5956 2728 6012
rect 2664 5952 2728 5956
rect 2744 6012 2808 6016
rect 2744 5956 2748 6012
rect 2748 5956 2804 6012
rect 2804 5956 2808 6012
rect 2744 5952 2808 5956
rect 2824 6012 2888 6016
rect 2824 5956 2828 6012
rect 2828 5956 2884 6012
rect 2884 5956 2888 6012
rect 2824 5952 2888 5956
rect 5847 6012 5911 6016
rect 5847 5956 5851 6012
rect 5851 5956 5907 6012
rect 5907 5956 5911 6012
rect 5847 5952 5911 5956
rect 5927 6012 5991 6016
rect 5927 5956 5931 6012
rect 5931 5956 5987 6012
rect 5987 5956 5991 6012
rect 5927 5952 5991 5956
rect 6007 6012 6071 6016
rect 6007 5956 6011 6012
rect 6011 5956 6067 6012
rect 6067 5956 6071 6012
rect 6007 5952 6071 5956
rect 6087 6012 6151 6016
rect 6087 5956 6091 6012
rect 6091 5956 6147 6012
rect 6147 5956 6151 6012
rect 6087 5952 6151 5956
rect 9111 6012 9175 6016
rect 9111 5956 9115 6012
rect 9115 5956 9171 6012
rect 9171 5956 9175 6012
rect 9111 5952 9175 5956
rect 9191 6012 9255 6016
rect 9191 5956 9195 6012
rect 9195 5956 9251 6012
rect 9251 5956 9255 6012
rect 9191 5952 9255 5956
rect 9271 6012 9335 6016
rect 9271 5956 9275 6012
rect 9275 5956 9331 6012
rect 9331 5956 9335 6012
rect 9271 5952 9335 5956
rect 9351 6012 9415 6016
rect 9351 5956 9355 6012
rect 9355 5956 9411 6012
rect 9411 5956 9415 6012
rect 9351 5952 9415 5956
rect 4215 5468 4279 5472
rect 4215 5412 4219 5468
rect 4219 5412 4275 5468
rect 4275 5412 4279 5468
rect 4215 5408 4279 5412
rect 4295 5468 4359 5472
rect 4295 5412 4299 5468
rect 4299 5412 4355 5468
rect 4355 5412 4359 5468
rect 4295 5408 4359 5412
rect 4375 5468 4439 5472
rect 4375 5412 4379 5468
rect 4379 5412 4435 5468
rect 4435 5412 4439 5468
rect 4375 5408 4439 5412
rect 4455 5468 4519 5472
rect 4455 5412 4459 5468
rect 4459 5412 4515 5468
rect 4515 5412 4519 5468
rect 4455 5408 4519 5412
rect 7479 5468 7543 5472
rect 7479 5412 7483 5468
rect 7483 5412 7539 5468
rect 7539 5412 7543 5468
rect 7479 5408 7543 5412
rect 7559 5468 7623 5472
rect 7559 5412 7563 5468
rect 7563 5412 7619 5468
rect 7619 5412 7623 5468
rect 7559 5408 7623 5412
rect 7639 5468 7703 5472
rect 7639 5412 7643 5468
rect 7643 5412 7699 5468
rect 7699 5412 7703 5468
rect 7639 5408 7703 5412
rect 7719 5468 7783 5472
rect 7719 5412 7723 5468
rect 7723 5412 7779 5468
rect 7779 5412 7783 5468
rect 7719 5408 7783 5412
rect 2584 4924 2648 4928
rect 2584 4868 2588 4924
rect 2588 4868 2644 4924
rect 2644 4868 2648 4924
rect 2584 4864 2648 4868
rect 2664 4924 2728 4928
rect 2664 4868 2668 4924
rect 2668 4868 2724 4924
rect 2724 4868 2728 4924
rect 2664 4864 2728 4868
rect 2744 4924 2808 4928
rect 2744 4868 2748 4924
rect 2748 4868 2804 4924
rect 2804 4868 2808 4924
rect 2744 4864 2808 4868
rect 2824 4924 2888 4928
rect 2824 4868 2828 4924
rect 2828 4868 2884 4924
rect 2884 4868 2888 4924
rect 2824 4864 2888 4868
rect 5847 4924 5911 4928
rect 5847 4868 5851 4924
rect 5851 4868 5907 4924
rect 5907 4868 5911 4924
rect 5847 4864 5911 4868
rect 5927 4924 5991 4928
rect 5927 4868 5931 4924
rect 5931 4868 5987 4924
rect 5987 4868 5991 4924
rect 5927 4864 5991 4868
rect 6007 4924 6071 4928
rect 6007 4868 6011 4924
rect 6011 4868 6067 4924
rect 6067 4868 6071 4924
rect 6007 4864 6071 4868
rect 6087 4924 6151 4928
rect 6087 4868 6091 4924
rect 6091 4868 6147 4924
rect 6147 4868 6151 4924
rect 6087 4864 6151 4868
rect 9111 4924 9175 4928
rect 9111 4868 9115 4924
rect 9115 4868 9171 4924
rect 9171 4868 9175 4924
rect 9111 4864 9175 4868
rect 9191 4924 9255 4928
rect 9191 4868 9195 4924
rect 9195 4868 9251 4924
rect 9251 4868 9255 4924
rect 9191 4864 9255 4868
rect 9271 4924 9335 4928
rect 9271 4868 9275 4924
rect 9275 4868 9331 4924
rect 9331 4868 9335 4924
rect 9271 4864 9335 4868
rect 9351 4924 9415 4928
rect 9351 4868 9355 4924
rect 9355 4868 9411 4924
rect 9411 4868 9415 4924
rect 9351 4864 9415 4868
rect 4215 4380 4279 4384
rect 4215 4324 4219 4380
rect 4219 4324 4275 4380
rect 4275 4324 4279 4380
rect 4215 4320 4279 4324
rect 4295 4380 4359 4384
rect 4295 4324 4299 4380
rect 4299 4324 4355 4380
rect 4355 4324 4359 4380
rect 4295 4320 4359 4324
rect 4375 4380 4439 4384
rect 4375 4324 4379 4380
rect 4379 4324 4435 4380
rect 4435 4324 4439 4380
rect 4375 4320 4439 4324
rect 4455 4380 4519 4384
rect 4455 4324 4459 4380
rect 4459 4324 4515 4380
rect 4515 4324 4519 4380
rect 4455 4320 4519 4324
rect 7479 4380 7543 4384
rect 7479 4324 7483 4380
rect 7483 4324 7539 4380
rect 7539 4324 7543 4380
rect 7479 4320 7543 4324
rect 7559 4380 7623 4384
rect 7559 4324 7563 4380
rect 7563 4324 7619 4380
rect 7619 4324 7623 4380
rect 7559 4320 7623 4324
rect 7639 4380 7703 4384
rect 7639 4324 7643 4380
rect 7643 4324 7699 4380
rect 7699 4324 7703 4380
rect 7639 4320 7703 4324
rect 7719 4380 7783 4384
rect 7719 4324 7723 4380
rect 7723 4324 7779 4380
rect 7779 4324 7783 4380
rect 7719 4320 7783 4324
rect 2584 3836 2648 3840
rect 2584 3780 2588 3836
rect 2588 3780 2644 3836
rect 2644 3780 2648 3836
rect 2584 3776 2648 3780
rect 2664 3836 2728 3840
rect 2664 3780 2668 3836
rect 2668 3780 2724 3836
rect 2724 3780 2728 3836
rect 2664 3776 2728 3780
rect 2744 3836 2808 3840
rect 2744 3780 2748 3836
rect 2748 3780 2804 3836
rect 2804 3780 2808 3836
rect 2744 3776 2808 3780
rect 2824 3836 2888 3840
rect 2824 3780 2828 3836
rect 2828 3780 2884 3836
rect 2884 3780 2888 3836
rect 2824 3776 2888 3780
rect 5847 3836 5911 3840
rect 5847 3780 5851 3836
rect 5851 3780 5907 3836
rect 5907 3780 5911 3836
rect 5847 3776 5911 3780
rect 5927 3836 5991 3840
rect 5927 3780 5931 3836
rect 5931 3780 5987 3836
rect 5987 3780 5991 3836
rect 5927 3776 5991 3780
rect 6007 3836 6071 3840
rect 6007 3780 6011 3836
rect 6011 3780 6067 3836
rect 6067 3780 6071 3836
rect 6007 3776 6071 3780
rect 6087 3836 6151 3840
rect 6087 3780 6091 3836
rect 6091 3780 6147 3836
rect 6147 3780 6151 3836
rect 6087 3776 6151 3780
rect 9111 3836 9175 3840
rect 9111 3780 9115 3836
rect 9115 3780 9171 3836
rect 9171 3780 9175 3836
rect 9111 3776 9175 3780
rect 9191 3836 9255 3840
rect 9191 3780 9195 3836
rect 9195 3780 9251 3836
rect 9251 3780 9255 3836
rect 9191 3776 9255 3780
rect 9271 3836 9335 3840
rect 9271 3780 9275 3836
rect 9275 3780 9331 3836
rect 9331 3780 9335 3836
rect 9271 3776 9335 3780
rect 9351 3836 9415 3840
rect 9351 3780 9355 3836
rect 9355 3780 9411 3836
rect 9411 3780 9415 3836
rect 9351 3776 9415 3780
rect 4215 3292 4279 3296
rect 4215 3236 4219 3292
rect 4219 3236 4275 3292
rect 4275 3236 4279 3292
rect 4215 3232 4279 3236
rect 4295 3292 4359 3296
rect 4295 3236 4299 3292
rect 4299 3236 4355 3292
rect 4355 3236 4359 3292
rect 4295 3232 4359 3236
rect 4375 3292 4439 3296
rect 4375 3236 4379 3292
rect 4379 3236 4435 3292
rect 4435 3236 4439 3292
rect 4375 3232 4439 3236
rect 4455 3292 4519 3296
rect 4455 3236 4459 3292
rect 4459 3236 4515 3292
rect 4515 3236 4519 3292
rect 4455 3232 4519 3236
rect 7479 3292 7543 3296
rect 7479 3236 7483 3292
rect 7483 3236 7539 3292
rect 7539 3236 7543 3292
rect 7479 3232 7543 3236
rect 7559 3292 7623 3296
rect 7559 3236 7563 3292
rect 7563 3236 7619 3292
rect 7619 3236 7623 3292
rect 7559 3232 7623 3236
rect 7639 3292 7703 3296
rect 7639 3236 7643 3292
rect 7643 3236 7699 3292
rect 7699 3236 7703 3292
rect 7639 3232 7703 3236
rect 7719 3292 7783 3296
rect 7719 3236 7723 3292
rect 7723 3236 7779 3292
rect 7779 3236 7783 3292
rect 7719 3232 7783 3236
rect 2584 2748 2648 2752
rect 2584 2692 2588 2748
rect 2588 2692 2644 2748
rect 2644 2692 2648 2748
rect 2584 2688 2648 2692
rect 2664 2748 2728 2752
rect 2664 2692 2668 2748
rect 2668 2692 2724 2748
rect 2724 2692 2728 2748
rect 2664 2688 2728 2692
rect 2744 2748 2808 2752
rect 2744 2692 2748 2748
rect 2748 2692 2804 2748
rect 2804 2692 2808 2748
rect 2744 2688 2808 2692
rect 2824 2748 2888 2752
rect 2824 2692 2828 2748
rect 2828 2692 2884 2748
rect 2884 2692 2888 2748
rect 2824 2688 2888 2692
rect 5847 2748 5911 2752
rect 5847 2692 5851 2748
rect 5851 2692 5907 2748
rect 5907 2692 5911 2748
rect 5847 2688 5911 2692
rect 5927 2748 5991 2752
rect 5927 2692 5931 2748
rect 5931 2692 5987 2748
rect 5987 2692 5991 2748
rect 5927 2688 5991 2692
rect 6007 2748 6071 2752
rect 6007 2692 6011 2748
rect 6011 2692 6067 2748
rect 6067 2692 6071 2748
rect 6007 2688 6071 2692
rect 6087 2748 6151 2752
rect 6087 2692 6091 2748
rect 6091 2692 6147 2748
rect 6147 2692 6151 2748
rect 6087 2688 6151 2692
rect 9111 2748 9175 2752
rect 9111 2692 9115 2748
rect 9115 2692 9171 2748
rect 9171 2692 9175 2748
rect 9111 2688 9175 2692
rect 9191 2748 9255 2752
rect 9191 2692 9195 2748
rect 9195 2692 9251 2748
rect 9251 2692 9255 2748
rect 9191 2688 9255 2692
rect 9271 2748 9335 2752
rect 9271 2692 9275 2748
rect 9275 2692 9331 2748
rect 9331 2692 9335 2748
rect 9271 2688 9335 2692
rect 9351 2748 9415 2752
rect 9351 2692 9355 2748
rect 9355 2692 9411 2748
rect 9411 2692 9415 2748
rect 9351 2688 9415 2692
rect 4215 2204 4279 2208
rect 4215 2148 4219 2204
rect 4219 2148 4275 2204
rect 4275 2148 4279 2204
rect 4215 2144 4279 2148
rect 4295 2204 4359 2208
rect 4295 2148 4299 2204
rect 4299 2148 4355 2204
rect 4355 2148 4359 2204
rect 4295 2144 4359 2148
rect 4375 2204 4439 2208
rect 4375 2148 4379 2204
rect 4379 2148 4435 2204
rect 4435 2148 4439 2204
rect 4375 2144 4439 2148
rect 4455 2204 4519 2208
rect 4455 2148 4459 2204
rect 4459 2148 4515 2204
rect 4515 2148 4519 2204
rect 4455 2144 4519 2148
rect 7479 2204 7543 2208
rect 7479 2148 7483 2204
rect 7483 2148 7539 2204
rect 7539 2148 7543 2204
rect 7479 2144 7543 2148
rect 7559 2204 7623 2208
rect 7559 2148 7563 2204
rect 7563 2148 7619 2204
rect 7619 2148 7623 2204
rect 7559 2144 7623 2148
rect 7639 2204 7703 2208
rect 7639 2148 7643 2204
rect 7643 2148 7699 2204
rect 7699 2148 7703 2204
rect 7639 2144 7703 2148
rect 7719 2204 7783 2208
rect 7719 2148 7723 2204
rect 7723 2148 7779 2204
rect 7779 2148 7783 2204
rect 7719 2144 7783 2148
<< metal4 >>
rect 2575 77824 2896 77840
rect 2575 77760 2584 77824
rect 2648 77760 2664 77824
rect 2728 77760 2744 77824
rect 2808 77760 2824 77824
rect 2888 77760 2896 77824
rect 2575 76736 2896 77760
rect 2575 76672 2584 76736
rect 2648 76672 2664 76736
rect 2728 76672 2744 76736
rect 2808 76672 2824 76736
rect 2888 76672 2896 76736
rect 2575 75648 2896 76672
rect 2575 75584 2584 75648
rect 2648 75584 2664 75648
rect 2728 75584 2744 75648
rect 2808 75584 2824 75648
rect 2888 75584 2896 75648
rect 2575 74560 2896 75584
rect 2575 74496 2584 74560
rect 2648 74496 2664 74560
rect 2728 74496 2744 74560
rect 2808 74496 2824 74560
rect 2888 74496 2896 74560
rect 2575 73472 2896 74496
rect 2575 73408 2584 73472
rect 2648 73408 2664 73472
rect 2728 73408 2744 73472
rect 2808 73408 2824 73472
rect 2888 73408 2896 73472
rect 2575 72384 2896 73408
rect 2575 72320 2584 72384
rect 2648 72320 2664 72384
rect 2728 72320 2744 72384
rect 2808 72320 2824 72384
rect 2888 72320 2896 72384
rect 2575 71296 2896 72320
rect 2575 71232 2584 71296
rect 2648 71232 2664 71296
rect 2728 71232 2744 71296
rect 2808 71232 2824 71296
rect 2888 71232 2896 71296
rect 2575 70208 2896 71232
rect 2575 70144 2584 70208
rect 2648 70144 2664 70208
rect 2728 70144 2744 70208
rect 2808 70144 2824 70208
rect 2888 70144 2896 70208
rect 2575 69120 2896 70144
rect 2575 69056 2584 69120
rect 2648 69056 2664 69120
rect 2728 69056 2744 69120
rect 2808 69056 2824 69120
rect 2888 69056 2896 69120
rect 1163 69052 1229 69053
rect 1163 68988 1164 69052
rect 1228 68988 1229 69052
rect 1163 68987 1229 68988
rect 1166 41173 1226 68987
rect 2575 68032 2896 69056
rect 2575 67968 2584 68032
rect 2648 67968 2664 68032
rect 2728 67968 2744 68032
rect 2808 67968 2824 68032
rect 2888 67968 2896 68032
rect 2575 66944 2896 67968
rect 2575 66880 2584 66944
rect 2648 66880 2664 66944
rect 2728 66880 2744 66944
rect 2808 66880 2824 66944
rect 2888 66880 2896 66944
rect 2575 65856 2896 66880
rect 2575 65792 2584 65856
rect 2648 65792 2664 65856
rect 2728 65792 2744 65856
rect 2808 65792 2824 65856
rect 2888 65792 2896 65856
rect 2575 64768 2896 65792
rect 2575 64704 2584 64768
rect 2648 64704 2664 64768
rect 2728 64704 2744 64768
rect 2808 64704 2824 64768
rect 2888 64704 2896 64768
rect 2575 63680 2896 64704
rect 2575 63616 2584 63680
rect 2648 63616 2664 63680
rect 2728 63616 2744 63680
rect 2808 63616 2824 63680
rect 2888 63616 2896 63680
rect 2575 62592 2896 63616
rect 2575 62528 2584 62592
rect 2648 62528 2664 62592
rect 2728 62528 2744 62592
rect 2808 62528 2824 62592
rect 2888 62528 2896 62592
rect 2575 61504 2896 62528
rect 2575 61440 2584 61504
rect 2648 61440 2664 61504
rect 2728 61440 2744 61504
rect 2808 61440 2824 61504
rect 2888 61440 2896 61504
rect 2575 60416 2896 61440
rect 2575 60352 2584 60416
rect 2648 60352 2664 60416
rect 2728 60352 2744 60416
rect 2808 60352 2824 60416
rect 2888 60352 2896 60416
rect 2575 59328 2896 60352
rect 2575 59264 2584 59328
rect 2648 59264 2664 59328
rect 2728 59264 2744 59328
rect 2808 59264 2824 59328
rect 2888 59264 2896 59328
rect 2575 58240 2896 59264
rect 2575 58176 2584 58240
rect 2648 58176 2664 58240
rect 2728 58176 2744 58240
rect 2808 58176 2824 58240
rect 2888 58176 2896 58240
rect 2267 57356 2333 57357
rect 2267 57292 2268 57356
rect 2332 57292 2333 57356
rect 2267 57291 2333 57292
rect 1899 54636 1965 54637
rect 1899 54572 1900 54636
rect 1964 54572 1965 54636
rect 1899 54571 1965 54572
rect 1902 50693 1962 54571
rect 2083 51100 2149 51101
rect 2083 51036 2084 51100
rect 2148 51036 2149 51100
rect 2083 51035 2149 51036
rect 1899 50692 1965 50693
rect 1899 50628 1900 50692
rect 1964 50628 1965 50692
rect 1899 50627 1965 50628
rect 2086 49061 2146 51035
rect 2270 50829 2330 57291
rect 2575 57152 2896 58176
rect 4207 77280 4527 77840
rect 4207 77216 4215 77280
rect 4279 77216 4295 77280
rect 4359 77216 4375 77280
rect 4439 77216 4455 77280
rect 4519 77216 4527 77280
rect 4207 76192 4527 77216
rect 4207 76128 4215 76192
rect 4279 76128 4295 76192
rect 4359 76128 4375 76192
rect 4439 76128 4455 76192
rect 4519 76128 4527 76192
rect 4207 75104 4527 76128
rect 4207 75040 4215 75104
rect 4279 75040 4295 75104
rect 4359 75040 4375 75104
rect 4439 75040 4455 75104
rect 4519 75040 4527 75104
rect 4207 74016 4527 75040
rect 4207 73952 4215 74016
rect 4279 73952 4295 74016
rect 4359 73952 4375 74016
rect 4439 73952 4455 74016
rect 4519 73952 4527 74016
rect 4207 72928 4527 73952
rect 4207 72864 4215 72928
rect 4279 72864 4295 72928
rect 4359 72864 4375 72928
rect 4439 72864 4455 72928
rect 4519 72864 4527 72928
rect 4207 71840 4527 72864
rect 4207 71776 4215 71840
rect 4279 71776 4295 71840
rect 4359 71776 4375 71840
rect 4439 71776 4455 71840
rect 4519 71776 4527 71840
rect 4207 70752 4527 71776
rect 4207 70688 4215 70752
rect 4279 70688 4295 70752
rect 4359 70688 4375 70752
rect 4439 70688 4455 70752
rect 4519 70688 4527 70752
rect 4207 69664 4527 70688
rect 4207 69600 4215 69664
rect 4279 69600 4295 69664
rect 4359 69600 4375 69664
rect 4439 69600 4455 69664
rect 4519 69600 4527 69664
rect 4207 68576 4527 69600
rect 4207 68512 4215 68576
rect 4279 68512 4295 68576
rect 4359 68512 4375 68576
rect 4439 68512 4455 68576
rect 4519 68512 4527 68576
rect 4207 67488 4527 68512
rect 4207 67424 4215 67488
rect 4279 67424 4295 67488
rect 4359 67424 4375 67488
rect 4439 67424 4455 67488
rect 4519 67424 4527 67488
rect 4207 66400 4527 67424
rect 4207 66336 4215 66400
rect 4279 66336 4295 66400
rect 4359 66336 4375 66400
rect 4439 66336 4455 66400
rect 4519 66336 4527 66400
rect 4207 65312 4527 66336
rect 4207 65248 4215 65312
rect 4279 65248 4295 65312
rect 4359 65248 4375 65312
rect 4439 65248 4455 65312
rect 4519 65248 4527 65312
rect 4207 64224 4527 65248
rect 4207 64160 4215 64224
rect 4279 64160 4295 64224
rect 4359 64160 4375 64224
rect 4439 64160 4455 64224
rect 4519 64160 4527 64224
rect 4207 63136 4527 64160
rect 4207 63072 4215 63136
rect 4279 63072 4295 63136
rect 4359 63072 4375 63136
rect 4439 63072 4455 63136
rect 4519 63072 4527 63136
rect 4207 62048 4527 63072
rect 4207 61984 4215 62048
rect 4279 61984 4295 62048
rect 4359 61984 4375 62048
rect 4439 61984 4455 62048
rect 4519 61984 4527 62048
rect 4207 60960 4527 61984
rect 4207 60896 4215 60960
rect 4279 60896 4295 60960
rect 4359 60896 4375 60960
rect 4439 60896 4455 60960
rect 4519 60896 4527 60960
rect 4207 59872 4527 60896
rect 4207 59808 4215 59872
rect 4279 59808 4295 59872
rect 4359 59808 4375 59872
rect 4439 59808 4455 59872
rect 4519 59808 4527 59872
rect 4207 58784 4527 59808
rect 4207 58720 4215 58784
rect 4279 58720 4295 58784
rect 4359 58720 4375 58784
rect 4439 58720 4455 58784
rect 4519 58720 4527 58784
rect 4207 57696 4527 58720
rect 4207 57632 4215 57696
rect 4279 57632 4295 57696
rect 4359 57632 4375 57696
rect 4439 57632 4455 57696
rect 4519 57632 4527 57696
rect 3187 57628 3253 57629
rect 3187 57564 3188 57628
rect 3252 57564 3253 57628
rect 3187 57563 3253 57564
rect 2575 57088 2584 57152
rect 2648 57088 2664 57152
rect 2728 57088 2744 57152
rect 2808 57088 2824 57152
rect 2888 57088 2896 57152
rect 2575 56064 2896 57088
rect 2575 56000 2584 56064
rect 2648 56000 2664 56064
rect 2728 56000 2744 56064
rect 2808 56000 2824 56064
rect 2888 56000 2896 56064
rect 2575 54976 2896 56000
rect 3190 55453 3250 57563
rect 4207 56608 4527 57632
rect 4207 56544 4215 56608
rect 4279 56544 4295 56608
rect 4359 56544 4375 56608
rect 4439 56544 4455 56608
rect 4519 56544 4527 56608
rect 3371 56268 3437 56269
rect 3371 56204 3372 56268
rect 3436 56204 3437 56268
rect 3371 56203 3437 56204
rect 3187 55452 3253 55453
rect 3187 55388 3188 55452
rect 3252 55388 3253 55452
rect 3187 55387 3253 55388
rect 2575 54912 2584 54976
rect 2648 54912 2664 54976
rect 2728 54912 2744 54976
rect 2808 54912 2824 54976
rect 2888 54912 2896 54976
rect 2575 53888 2896 54912
rect 2575 53824 2584 53888
rect 2648 53824 2664 53888
rect 2728 53824 2744 53888
rect 2808 53824 2824 53888
rect 2888 53824 2896 53888
rect 2575 52800 2896 53824
rect 2575 52736 2584 52800
rect 2648 52736 2664 52800
rect 2728 52736 2744 52800
rect 2808 52736 2824 52800
rect 2888 52736 2896 52800
rect 2575 51712 2896 52736
rect 2575 51648 2584 51712
rect 2648 51648 2664 51712
rect 2728 51648 2744 51712
rect 2808 51648 2824 51712
rect 2888 51648 2896 51712
rect 2267 50828 2333 50829
rect 2267 50764 2268 50828
rect 2332 50764 2333 50828
rect 2267 50763 2333 50764
rect 2575 50624 2896 51648
rect 3003 50828 3069 50829
rect 3003 50764 3004 50828
rect 3068 50764 3069 50828
rect 3003 50763 3069 50764
rect 2575 50560 2584 50624
rect 2648 50560 2664 50624
rect 2728 50560 2744 50624
rect 2808 50560 2824 50624
rect 2888 50560 2896 50624
rect 2575 49536 2896 50560
rect 2575 49472 2584 49536
rect 2648 49472 2664 49536
rect 2728 49472 2744 49536
rect 2808 49472 2824 49536
rect 2888 49472 2896 49536
rect 2083 49060 2149 49061
rect 2083 48996 2084 49060
rect 2148 48996 2149 49060
rect 2083 48995 2149 48996
rect 2575 48448 2896 49472
rect 2575 48384 2584 48448
rect 2648 48384 2664 48448
rect 2728 48384 2744 48448
rect 2808 48384 2824 48448
rect 2888 48384 2896 48448
rect 2267 48244 2333 48245
rect 2267 48180 2268 48244
rect 2332 48180 2333 48244
rect 2267 48179 2333 48180
rect 2083 45116 2149 45117
rect 2083 45052 2084 45116
rect 2148 45052 2149 45116
rect 2083 45051 2149 45052
rect 2086 42125 2146 45051
rect 2270 43485 2330 48179
rect 2575 47360 2896 48384
rect 2575 47296 2584 47360
rect 2648 47296 2664 47360
rect 2728 47296 2744 47360
rect 2808 47296 2824 47360
rect 2888 47296 2896 47360
rect 2575 46272 2896 47296
rect 2575 46208 2584 46272
rect 2648 46208 2664 46272
rect 2728 46208 2744 46272
rect 2808 46208 2824 46272
rect 2888 46208 2896 46272
rect 2575 45184 2896 46208
rect 3006 46069 3066 50763
rect 3190 50557 3250 55387
rect 3374 50829 3434 56203
rect 4207 55520 4527 56544
rect 4207 55456 4215 55520
rect 4279 55456 4295 55520
rect 4359 55456 4375 55520
rect 4439 55456 4455 55520
rect 4519 55456 4527 55520
rect 4207 54432 4527 55456
rect 4207 54368 4215 54432
rect 4279 54368 4295 54432
rect 4359 54368 4375 54432
rect 4439 54368 4455 54432
rect 4519 54368 4527 54432
rect 4207 53344 4527 54368
rect 4207 53280 4215 53344
rect 4279 53280 4295 53344
rect 4359 53280 4375 53344
rect 4439 53280 4455 53344
rect 4519 53280 4527 53344
rect 4207 52256 4527 53280
rect 4207 52192 4215 52256
rect 4279 52192 4295 52256
rect 4359 52192 4375 52256
rect 4439 52192 4455 52256
rect 4519 52192 4527 52256
rect 3923 51236 3989 51237
rect 3923 51172 3924 51236
rect 3988 51172 3989 51236
rect 3923 51171 3989 51172
rect 3739 51100 3805 51101
rect 3739 51036 3740 51100
rect 3804 51036 3805 51100
rect 3739 51035 3805 51036
rect 3371 50828 3437 50829
rect 3371 50764 3372 50828
rect 3436 50764 3437 50828
rect 3371 50763 3437 50764
rect 3187 50556 3253 50557
rect 3187 50492 3188 50556
rect 3252 50492 3253 50556
rect 3187 50491 3253 50492
rect 3742 49605 3802 51035
rect 3926 49877 3986 51171
rect 4207 51168 4527 52192
rect 4207 51104 4215 51168
rect 4279 51104 4295 51168
rect 4359 51104 4375 51168
rect 4439 51104 4455 51168
rect 4519 51104 4527 51168
rect 4207 50080 4527 51104
rect 4207 50016 4215 50080
rect 4279 50016 4295 50080
rect 4359 50016 4375 50080
rect 4439 50016 4455 50080
rect 4519 50016 4527 50080
rect 3923 49876 3989 49877
rect 3923 49812 3924 49876
rect 3988 49812 3989 49876
rect 3923 49811 3989 49812
rect 3739 49604 3805 49605
rect 3739 49540 3740 49604
rect 3804 49540 3805 49604
rect 3739 49539 3805 49540
rect 4207 48992 4527 50016
rect 5839 77824 6159 77840
rect 5839 77760 5847 77824
rect 5911 77760 5927 77824
rect 5991 77760 6007 77824
rect 6071 77760 6087 77824
rect 6151 77760 6159 77824
rect 5839 76736 6159 77760
rect 5839 76672 5847 76736
rect 5911 76672 5927 76736
rect 5991 76672 6007 76736
rect 6071 76672 6087 76736
rect 6151 76672 6159 76736
rect 5839 75648 6159 76672
rect 5839 75584 5847 75648
rect 5911 75584 5927 75648
rect 5991 75584 6007 75648
rect 6071 75584 6087 75648
rect 6151 75584 6159 75648
rect 5839 74560 6159 75584
rect 5839 74496 5847 74560
rect 5911 74496 5927 74560
rect 5991 74496 6007 74560
rect 6071 74496 6087 74560
rect 6151 74496 6159 74560
rect 5839 73472 6159 74496
rect 5839 73408 5847 73472
rect 5911 73408 5927 73472
rect 5991 73408 6007 73472
rect 6071 73408 6087 73472
rect 6151 73408 6159 73472
rect 5839 72384 6159 73408
rect 5839 72320 5847 72384
rect 5911 72320 5927 72384
rect 5991 72320 6007 72384
rect 6071 72320 6087 72384
rect 6151 72320 6159 72384
rect 5839 71296 6159 72320
rect 5839 71232 5847 71296
rect 5911 71232 5927 71296
rect 5991 71232 6007 71296
rect 6071 71232 6087 71296
rect 6151 71232 6159 71296
rect 5839 70208 6159 71232
rect 5839 70144 5847 70208
rect 5911 70144 5927 70208
rect 5991 70144 6007 70208
rect 6071 70144 6087 70208
rect 6151 70144 6159 70208
rect 5839 69120 6159 70144
rect 5839 69056 5847 69120
rect 5911 69056 5927 69120
rect 5991 69056 6007 69120
rect 6071 69056 6087 69120
rect 6151 69056 6159 69120
rect 5839 68032 6159 69056
rect 5839 67968 5847 68032
rect 5911 67968 5927 68032
rect 5991 67968 6007 68032
rect 6071 67968 6087 68032
rect 6151 67968 6159 68032
rect 5839 66944 6159 67968
rect 5839 66880 5847 66944
rect 5911 66880 5927 66944
rect 5991 66880 6007 66944
rect 6071 66880 6087 66944
rect 6151 66880 6159 66944
rect 5839 65856 6159 66880
rect 5839 65792 5847 65856
rect 5911 65792 5927 65856
rect 5991 65792 6007 65856
rect 6071 65792 6087 65856
rect 6151 65792 6159 65856
rect 5839 64768 6159 65792
rect 5839 64704 5847 64768
rect 5911 64704 5927 64768
rect 5991 64704 6007 64768
rect 6071 64704 6087 64768
rect 6151 64704 6159 64768
rect 5839 63680 6159 64704
rect 5839 63616 5847 63680
rect 5911 63616 5927 63680
rect 5991 63616 6007 63680
rect 6071 63616 6087 63680
rect 6151 63616 6159 63680
rect 5839 62592 6159 63616
rect 5839 62528 5847 62592
rect 5911 62528 5927 62592
rect 5991 62528 6007 62592
rect 6071 62528 6087 62592
rect 6151 62528 6159 62592
rect 5839 61504 6159 62528
rect 5839 61440 5847 61504
rect 5911 61440 5927 61504
rect 5991 61440 6007 61504
rect 6071 61440 6087 61504
rect 6151 61440 6159 61504
rect 5839 60416 6159 61440
rect 5839 60352 5847 60416
rect 5911 60352 5927 60416
rect 5991 60352 6007 60416
rect 6071 60352 6087 60416
rect 6151 60352 6159 60416
rect 5839 59328 6159 60352
rect 5839 59264 5847 59328
rect 5911 59264 5927 59328
rect 5991 59264 6007 59328
rect 6071 59264 6087 59328
rect 6151 59264 6159 59328
rect 5839 58240 6159 59264
rect 5839 58176 5847 58240
rect 5911 58176 5927 58240
rect 5991 58176 6007 58240
rect 6071 58176 6087 58240
rect 6151 58176 6159 58240
rect 5839 57152 6159 58176
rect 5839 57088 5847 57152
rect 5911 57088 5927 57152
rect 5991 57088 6007 57152
rect 6071 57088 6087 57152
rect 6151 57088 6159 57152
rect 5839 56064 6159 57088
rect 5839 56000 5847 56064
rect 5911 56000 5927 56064
rect 5991 56000 6007 56064
rect 6071 56000 6087 56064
rect 6151 56000 6159 56064
rect 5839 54976 6159 56000
rect 5839 54912 5847 54976
rect 5911 54912 5927 54976
rect 5991 54912 6007 54976
rect 6071 54912 6087 54976
rect 6151 54912 6159 54976
rect 5839 53888 6159 54912
rect 5839 53824 5847 53888
rect 5911 53824 5927 53888
rect 5991 53824 6007 53888
rect 6071 53824 6087 53888
rect 6151 53824 6159 53888
rect 5839 52800 6159 53824
rect 5839 52736 5847 52800
rect 5911 52736 5927 52800
rect 5991 52736 6007 52800
rect 6071 52736 6087 52800
rect 6151 52736 6159 52800
rect 5839 51712 6159 52736
rect 5839 51648 5847 51712
rect 5911 51648 5927 51712
rect 5991 51648 6007 51712
rect 6071 51648 6087 51712
rect 6151 51648 6159 51712
rect 5839 50624 6159 51648
rect 7471 77280 7791 77840
rect 7471 77216 7479 77280
rect 7543 77216 7559 77280
rect 7623 77216 7639 77280
rect 7703 77216 7719 77280
rect 7783 77216 7791 77280
rect 7471 76192 7791 77216
rect 7471 76128 7479 76192
rect 7543 76128 7559 76192
rect 7623 76128 7639 76192
rect 7703 76128 7719 76192
rect 7783 76128 7791 76192
rect 7471 75104 7791 76128
rect 7471 75040 7479 75104
rect 7543 75040 7559 75104
rect 7623 75040 7639 75104
rect 7703 75040 7719 75104
rect 7783 75040 7791 75104
rect 7471 74016 7791 75040
rect 7471 73952 7479 74016
rect 7543 73952 7559 74016
rect 7623 73952 7639 74016
rect 7703 73952 7719 74016
rect 7783 73952 7791 74016
rect 7471 72928 7791 73952
rect 7471 72864 7479 72928
rect 7543 72864 7559 72928
rect 7623 72864 7639 72928
rect 7703 72864 7719 72928
rect 7783 72864 7791 72928
rect 7471 71840 7791 72864
rect 7471 71776 7479 71840
rect 7543 71776 7559 71840
rect 7623 71776 7639 71840
rect 7703 71776 7719 71840
rect 7783 71776 7791 71840
rect 7471 70752 7791 71776
rect 7471 70688 7479 70752
rect 7543 70688 7559 70752
rect 7623 70688 7639 70752
rect 7703 70688 7719 70752
rect 7783 70688 7791 70752
rect 7471 69664 7791 70688
rect 7471 69600 7479 69664
rect 7543 69600 7559 69664
rect 7623 69600 7639 69664
rect 7703 69600 7719 69664
rect 7783 69600 7791 69664
rect 7471 68576 7791 69600
rect 7471 68512 7479 68576
rect 7543 68512 7559 68576
rect 7623 68512 7639 68576
rect 7703 68512 7719 68576
rect 7783 68512 7791 68576
rect 7471 67488 7791 68512
rect 7471 67424 7479 67488
rect 7543 67424 7559 67488
rect 7623 67424 7639 67488
rect 7703 67424 7719 67488
rect 7783 67424 7791 67488
rect 7471 66400 7791 67424
rect 7471 66336 7479 66400
rect 7543 66336 7559 66400
rect 7623 66336 7639 66400
rect 7703 66336 7719 66400
rect 7783 66336 7791 66400
rect 7471 65312 7791 66336
rect 7471 65248 7479 65312
rect 7543 65248 7559 65312
rect 7623 65248 7639 65312
rect 7703 65248 7719 65312
rect 7783 65248 7791 65312
rect 7471 64224 7791 65248
rect 7471 64160 7479 64224
rect 7543 64160 7559 64224
rect 7623 64160 7639 64224
rect 7703 64160 7719 64224
rect 7783 64160 7791 64224
rect 7471 63136 7791 64160
rect 7471 63072 7479 63136
rect 7543 63072 7559 63136
rect 7623 63072 7639 63136
rect 7703 63072 7719 63136
rect 7783 63072 7791 63136
rect 7471 62048 7791 63072
rect 7471 61984 7479 62048
rect 7543 61984 7559 62048
rect 7623 61984 7639 62048
rect 7703 61984 7719 62048
rect 7783 61984 7791 62048
rect 7471 60960 7791 61984
rect 7471 60896 7479 60960
rect 7543 60896 7559 60960
rect 7623 60896 7639 60960
rect 7703 60896 7719 60960
rect 7783 60896 7791 60960
rect 7471 59872 7791 60896
rect 7471 59808 7479 59872
rect 7543 59808 7559 59872
rect 7623 59808 7639 59872
rect 7703 59808 7719 59872
rect 7783 59808 7791 59872
rect 7471 58784 7791 59808
rect 7471 58720 7479 58784
rect 7543 58720 7559 58784
rect 7623 58720 7639 58784
rect 7703 58720 7719 58784
rect 7783 58720 7791 58784
rect 7471 57696 7791 58720
rect 7471 57632 7479 57696
rect 7543 57632 7559 57696
rect 7623 57632 7639 57696
rect 7703 57632 7719 57696
rect 7783 57632 7791 57696
rect 7471 56608 7791 57632
rect 7471 56544 7479 56608
rect 7543 56544 7559 56608
rect 7623 56544 7639 56608
rect 7703 56544 7719 56608
rect 7783 56544 7791 56608
rect 7471 55520 7791 56544
rect 7471 55456 7479 55520
rect 7543 55456 7559 55520
rect 7623 55456 7639 55520
rect 7703 55456 7719 55520
rect 7783 55456 7791 55520
rect 7471 54432 7791 55456
rect 7471 54368 7479 54432
rect 7543 54368 7559 54432
rect 7623 54368 7639 54432
rect 7703 54368 7719 54432
rect 7783 54368 7791 54432
rect 7471 53344 7791 54368
rect 7471 53280 7479 53344
rect 7543 53280 7559 53344
rect 7623 53280 7639 53344
rect 7703 53280 7719 53344
rect 7783 53280 7791 53344
rect 7471 52256 7791 53280
rect 7471 52192 7479 52256
rect 7543 52192 7559 52256
rect 7623 52192 7639 52256
rect 7703 52192 7719 52256
rect 7783 52192 7791 52256
rect 7471 51168 7791 52192
rect 7471 51104 7479 51168
rect 7543 51104 7559 51168
rect 7623 51104 7639 51168
rect 7703 51104 7719 51168
rect 7783 51104 7791 51168
rect 6315 50964 6381 50965
rect 6315 50900 6316 50964
rect 6380 50900 6381 50964
rect 6315 50899 6381 50900
rect 5839 50560 5847 50624
rect 5911 50560 5927 50624
rect 5991 50560 6007 50624
rect 6071 50560 6087 50624
rect 6151 50560 6159 50624
rect 4659 49604 4725 49605
rect 4659 49540 4660 49604
rect 4724 49540 4725 49604
rect 4659 49539 4725 49540
rect 4207 48928 4215 48992
rect 4279 48928 4295 48992
rect 4359 48928 4375 48992
rect 4439 48928 4455 48992
rect 4519 48928 4527 48992
rect 4207 47904 4527 48928
rect 4207 47840 4215 47904
rect 4279 47840 4295 47904
rect 4359 47840 4375 47904
rect 4439 47840 4455 47904
rect 4519 47840 4527 47904
rect 4207 46816 4527 47840
rect 4207 46752 4215 46816
rect 4279 46752 4295 46816
rect 4359 46752 4375 46816
rect 4439 46752 4455 46816
rect 4519 46752 4527 46816
rect 3187 46748 3253 46749
rect 3187 46684 3188 46748
rect 3252 46684 3253 46748
rect 3187 46683 3253 46684
rect 3003 46068 3069 46069
rect 3003 46004 3004 46068
rect 3068 46004 3069 46068
rect 3003 46003 3069 46004
rect 2575 45120 2584 45184
rect 2648 45120 2664 45184
rect 2728 45120 2744 45184
rect 2808 45120 2824 45184
rect 2888 45120 2896 45184
rect 2575 44096 2896 45120
rect 3003 45116 3069 45117
rect 3003 45052 3004 45116
rect 3068 45052 3069 45116
rect 3003 45051 3069 45052
rect 2575 44032 2584 44096
rect 2648 44032 2664 44096
rect 2728 44032 2744 44096
rect 2808 44032 2824 44096
rect 2888 44032 2896 44096
rect 2267 43484 2333 43485
rect 2267 43420 2268 43484
rect 2332 43420 2333 43484
rect 2267 43419 2333 43420
rect 2575 43008 2896 44032
rect 2575 42944 2584 43008
rect 2648 42944 2664 43008
rect 2728 42944 2744 43008
rect 2808 42944 2824 43008
rect 2888 42944 2896 43008
rect 2083 42124 2149 42125
rect 2083 42060 2084 42124
rect 2148 42060 2149 42124
rect 2083 42059 2149 42060
rect 2575 41920 2896 42944
rect 2575 41856 2584 41920
rect 2648 41856 2664 41920
rect 2728 41856 2744 41920
rect 2808 41856 2824 41920
rect 2888 41856 2896 41920
rect 2267 41308 2333 41309
rect 2267 41244 2268 41308
rect 2332 41244 2333 41308
rect 2267 41243 2333 41244
rect 1163 41172 1229 41173
rect 1163 41108 1164 41172
rect 1228 41108 1229 41172
rect 1163 41107 1229 41108
rect 2083 38724 2149 38725
rect 2083 38660 2084 38724
rect 2148 38660 2149 38724
rect 2083 38659 2149 38660
rect 1531 36140 1597 36141
rect 1531 36076 1532 36140
rect 1596 36076 1597 36140
rect 1531 36075 1597 36076
rect 1534 32061 1594 36075
rect 2086 32469 2146 38659
rect 2270 32605 2330 41243
rect 2575 40832 2896 41856
rect 2575 40768 2584 40832
rect 2648 40768 2664 40832
rect 2728 40768 2744 40832
rect 2808 40768 2824 40832
rect 2888 40768 2896 40832
rect 2575 39744 2896 40768
rect 2575 39680 2584 39744
rect 2648 39680 2664 39744
rect 2728 39680 2744 39744
rect 2808 39680 2824 39744
rect 2888 39680 2896 39744
rect 2575 38656 2896 39680
rect 3006 38725 3066 45051
rect 3190 43349 3250 46683
rect 3923 46476 3989 46477
rect 3923 46412 3924 46476
rect 3988 46412 3989 46476
rect 3923 46411 3989 46412
rect 3187 43348 3253 43349
rect 3187 43284 3188 43348
rect 3252 43284 3253 43348
rect 3187 43283 3253 43284
rect 3926 38861 3986 46411
rect 4207 45728 4527 46752
rect 4207 45664 4215 45728
rect 4279 45664 4295 45728
rect 4359 45664 4375 45728
rect 4439 45664 4455 45728
rect 4519 45664 4527 45728
rect 4207 44640 4527 45664
rect 4207 44576 4215 44640
rect 4279 44576 4295 44640
rect 4359 44576 4375 44640
rect 4439 44576 4455 44640
rect 4519 44576 4527 44640
rect 4207 43552 4527 44576
rect 4207 43488 4215 43552
rect 4279 43488 4295 43552
rect 4359 43488 4375 43552
rect 4439 43488 4455 43552
rect 4519 43488 4527 43552
rect 4207 42464 4527 43488
rect 4662 43349 4722 49539
rect 5839 49536 6159 50560
rect 5839 49472 5847 49536
rect 5911 49472 5927 49536
rect 5991 49472 6007 49536
rect 6071 49472 6087 49536
rect 6151 49472 6159 49536
rect 5395 49060 5461 49061
rect 5395 48996 5396 49060
rect 5460 48996 5461 49060
rect 5395 48995 5461 48996
rect 5398 48517 5458 48995
rect 5579 48924 5645 48925
rect 5579 48860 5580 48924
rect 5644 48860 5645 48924
rect 5579 48859 5645 48860
rect 5395 48516 5461 48517
rect 5395 48452 5396 48516
rect 5460 48452 5461 48516
rect 5395 48451 5461 48452
rect 5582 48381 5642 48859
rect 5839 48448 6159 49472
rect 5839 48384 5847 48448
rect 5911 48384 5927 48448
rect 5991 48384 6007 48448
rect 6071 48384 6087 48448
rect 6151 48384 6159 48448
rect 5579 48380 5645 48381
rect 5579 48316 5580 48380
rect 5644 48316 5645 48380
rect 5579 48315 5645 48316
rect 4843 47836 4909 47837
rect 4843 47772 4844 47836
rect 4908 47772 4909 47836
rect 4843 47771 4909 47772
rect 4659 43348 4725 43349
rect 4659 43284 4660 43348
rect 4724 43284 4725 43348
rect 4659 43283 4725 43284
rect 4207 42400 4215 42464
rect 4279 42400 4295 42464
rect 4359 42400 4375 42464
rect 4439 42400 4455 42464
rect 4519 42400 4527 42464
rect 4207 41376 4527 42400
rect 4846 42261 4906 47771
rect 5839 47360 6159 48384
rect 5839 47296 5847 47360
rect 5911 47296 5927 47360
rect 5991 47296 6007 47360
rect 6071 47296 6087 47360
rect 6151 47296 6159 47360
rect 5839 46272 6159 47296
rect 5839 46208 5847 46272
rect 5911 46208 5927 46272
rect 5991 46208 6007 46272
rect 6071 46208 6087 46272
rect 6151 46208 6159 46272
rect 5027 46204 5093 46205
rect 5027 46140 5028 46204
rect 5092 46140 5093 46204
rect 5027 46139 5093 46140
rect 4843 42260 4909 42261
rect 4843 42196 4844 42260
rect 4908 42196 4909 42260
rect 4843 42195 4909 42196
rect 5030 41989 5090 46139
rect 5839 45184 6159 46208
rect 5839 45120 5847 45184
rect 5911 45120 5927 45184
rect 5991 45120 6007 45184
rect 6071 45120 6087 45184
rect 6151 45120 6159 45184
rect 5839 44096 6159 45120
rect 5839 44032 5847 44096
rect 5911 44032 5927 44096
rect 5991 44032 6007 44096
rect 6071 44032 6087 44096
rect 6151 44032 6159 44096
rect 5839 43008 6159 44032
rect 5839 42944 5847 43008
rect 5911 42944 5927 43008
rect 5991 42944 6007 43008
rect 6071 42944 6087 43008
rect 6151 42944 6159 43008
rect 5027 41988 5093 41989
rect 5027 41924 5028 41988
rect 5092 41924 5093 41988
rect 5027 41923 5093 41924
rect 5839 41920 6159 42944
rect 5839 41856 5847 41920
rect 5911 41856 5927 41920
rect 5991 41856 6007 41920
rect 6071 41856 6087 41920
rect 6151 41856 6159 41920
rect 5395 41716 5461 41717
rect 5395 41652 5396 41716
rect 5460 41652 5461 41716
rect 5395 41651 5461 41652
rect 5211 41580 5277 41581
rect 5211 41516 5212 41580
rect 5276 41516 5277 41580
rect 5211 41515 5277 41516
rect 4207 41312 4215 41376
rect 4279 41312 4295 41376
rect 4359 41312 4375 41376
rect 4439 41312 4455 41376
rect 4519 41312 4527 41376
rect 4207 40288 4527 41312
rect 4207 40224 4215 40288
rect 4279 40224 4295 40288
rect 4359 40224 4375 40288
rect 4439 40224 4455 40288
rect 4519 40224 4527 40288
rect 4207 39200 4527 40224
rect 5214 39813 5274 41515
rect 5211 39812 5277 39813
rect 5211 39748 5212 39812
rect 5276 39748 5277 39812
rect 5211 39747 5277 39748
rect 5398 39541 5458 41651
rect 5839 40832 6159 41856
rect 6318 41581 6378 50899
rect 7471 50080 7791 51104
rect 7471 50016 7479 50080
rect 7543 50016 7559 50080
rect 7623 50016 7639 50080
rect 7703 50016 7719 50080
rect 7783 50016 7791 50080
rect 6499 49740 6565 49741
rect 6499 49676 6500 49740
rect 6564 49676 6565 49740
rect 6499 49675 6565 49676
rect 6315 41580 6381 41581
rect 6315 41516 6316 41580
rect 6380 41516 6381 41580
rect 6315 41515 6381 41516
rect 6502 41309 6562 49675
rect 7471 48992 7791 50016
rect 7471 48928 7479 48992
rect 7543 48928 7559 48992
rect 7623 48928 7639 48992
rect 7703 48928 7719 48992
rect 7783 48928 7791 48992
rect 7471 47904 7791 48928
rect 7471 47840 7479 47904
rect 7543 47840 7559 47904
rect 7623 47840 7639 47904
rect 7703 47840 7719 47904
rect 7783 47840 7791 47904
rect 7471 46816 7791 47840
rect 7471 46752 7479 46816
rect 7543 46752 7559 46816
rect 7623 46752 7639 46816
rect 7703 46752 7719 46816
rect 7783 46752 7791 46816
rect 7471 45728 7791 46752
rect 7471 45664 7479 45728
rect 7543 45664 7559 45728
rect 7623 45664 7639 45728
rect 7703 45664 7719 45728
rect 7783 45664 7791 45728
rect 7471 44640 7791 45664
rect 7471 44576 7479 44640
rect 7543 44576 7559 44640
rect 7623 44576 7639 44640
rect 7703 44576 7719 44640
rect 7783 44576 7791 44640
rect 7471 43552 7791 44576
rect 7471 43488 7479 43552
rect 7543 43488 7559 43552
rect 7623 43488 7639 43552
rect 7703 43488 7719 43552
rect 7783 43488 7791 43552
rect 7471 42464 7791 43488
rect 7471 42400 7479 42464
rect 7543 42400 7559 42464
rect 7623 42400 7639 42464
rect 7703 42400 7719 42464
rect 7783 42400 7791 42464
rect 7471 41376 7791 42400
rect 7471 41312 7479 41376
rect 7543 41312 7559 41376
rect 7623 41312 7639 41376
rect 7703 41312 7719 41376
rect 7783 41312 7791 41376
rect 6499 41308 6565 41309
rect 6499 41244 6500 41308
rect 6564 41244 6565 41308
rect 6499 41243 6565 41244
rect 5839 40768 5847 40832
rect 5911 40768 5927 40832
rect 5991 40768 6007 40832
rect 6071 40768 6087 40832
rect 6151 40768 6159 40832
rect 5839 39744 6159 40768
rect 5839 39680 5847 39744
rect 5911 39680 5927 39744
rect 5991 39680 6007 39744
rect 6071 39680 6087 39744
rect 6151 39680 6159 39744
rect 5395 39540 5461 39541
rect 5395 39476 5396 39540
rect 5460 39476 5461 39540
rect 5395 39475 5461 39476
rect 4207 39136 4215 39200
rect 4279 39136 4295 39200
rect 4359 39136 4375 39200
rect 4439 39136 4455 39200
rect 4519 39136 4527 39200
rect 3923 38860 3989 38861
rect 3923 38796 3924 38860
rect 3988 38796 3989 38860
rect 3923 38795 3989 38796
rect 3003 38724 3069 38725
rect 3003 38660 3004 38724
rect 3068 38660 3069 38724
rect 3003 38659 3069 38660
rect 2575 38592 2584 38656
rect 2648 38592 2664 38656
rect 2728 38592 2744 38656
rect 2808 38592 2824 38656
rect 2888 38592 2896 38656
rect 2575 37568 2896 38592
rect 2575 37504 2584 37568
rect 2648 37504 2664 37568
rect 2728 37504 2744 37568
rect 2808 37504 2824 37568
rect 2888 37504 2896 37568
rect 2575 36480 2896 37504
rect 4207 38112 4527 39136
rect 4207 38048 4215 38112
rect 4279 38048 4295 38112
rect 4359 38048 4375 38112
rect 4439 38048 4455 38112
rect 4519 38048 4527 38112
rect 3739 37364 3805 37365
rect 3739 37300 3740 37364
rect 3804 37300 3805 37364
rect 3739 37299 3805 37300
rect 3003 37228 3069 37229
rect 3003 37164 3004 37228
rect 3068 37164 3069 37228
rect 3003 37163 3069 37164
rect 2575 36416 2584 36480
rect 2648 36416 2664 36480
rect 2728 36416 2744 36480
rect 2808 36416 2824 36480
rect 2888 36416 2896 36480
rect 2575 35392 2896 36416
rect 2575 35328 2584 35392
rect 2648 35328 2664 35392
rect 2728 35328 2744 35392
rect 2808 35328 2824 35392
rect 2888 35328 2896 35392
rect 2575 34304 2896 35328
rect 2575 34240 2584 34304
rect 2648 34240 2664 34304
rect 2728 34240 2744 34304
rect 2808 34240 2824 34304
rect 2888 34240 2896 34304
rect 2575 33216 2896 34240
rect 3006 33829 3066 37163
rect 3555 36684 3621 36685
rect 3555 36620 3556 36684
rect 3620 36620 3621 36684
rect 3555 36619 3621 36620
rect 3003 33828 3069 33829
rect 3003 33764 3004 33828
rect 3068 33764 3069 33828
rect 3003 33763 3069 33764
rect 2575 33152 2584 33216
rect 2648 33152 2664 33216
rect 2728 33152 2744 33216
rect 2808 33152 2824 33216
rect 2888 33152 2896 33216
rect 2267 32604 2333 32605
rect 2267 32540 2268 32604
rect 2332 32540 2333 32604
rect 2267 32539 2333 32540
rect 2083 32468 2149 32469
rect 2083 32404 2084 32468
rect 2148 32404 2149 32468
rect 2083 32403 2149 32404
rect 2575 32128 2896 33152
rect 2575 32064 2584 32128
rect 2648 32064 2664 32128
rect 2728 32064 2744 32128
rect 2808 32064 2824 32128
rect 2888 32064 2896 32128
rect 1531 32060 1597 32061
rect 1531 31996 1532 32060
rect 1596 31996 1597 32060
rect 1531 31995 1597 31996
rect 1715 31788 1781 31789
rect 1715 31724 1716 31788
rect 1780 31724 1781 31788
rect 1715 31723 1781 31724
rect 1718 29205 1778 31723
rect 2575 31040 2896 32064
rect 3558 31653 3618 36619
rect 3742 35461 3802 37299
rect 4207 37024 4527 38048
rect 4207 36960 4215 37024
rect 4279 36960 4295 37024
rect 4359 36960 4375 37024
rect 4439 36960 4455 37024
rect 4519 36960 4527 37024
rect 4207 35936 4527 36960
rect 4207 35872 4215 35936
rect 4279 35872 4295 35936
rect 4359 35872 4375 35936
rect 4439 35872 4455 35936
rect 4519 35872 4527 35936
rect 3739 35460 3805 35461
rect 3739 35396 3740 35460
rect 3804 35396 3805 35460
rect 3739 35395 3805 35396
rect 4207 34848 4527 35872
rect 4207 34784 4215 34848
rect 4279 34784 4295 34848
rect 4359 34784 4375 34848
rect 4439 34784 4455 34848
rect 4519 34784 4527 34848
rect 4207 33760 4527 34784
rect 4207 33696 4215 33760
rect 4279 33696 4295 33760
rect 4359 33696 4375 33760
rect 4439 33696 4455 33760
rect 4519 33696 4527 33760
rect 4207 32672 4527 33696
rect 4207 32608 4215 32672
rect 4279 32608 4295 32672
rect 4359 32608 4375 32672
rect 4439 32608 4455 32672
rect 4519 32608 4527 32672
rect 3555 31652 3621 31653
rect 3555 31588 3556 31652
rect 3620 31588 3621 31652
rect 3555 31587 3621 31588
rect 2575 30976 2584 31040
rect 2648 30976 2664 31040
rect 2728 30976 2744 31040
rect 2808 30976 2824 31040
rect 2888 30976 2896 31040
rect 2575 29952 2896 30976
rect 2575 29888 2584 29952
rect 2648 29888 2664 29952
rect 2728 29888 2744 29952
rect 2808 29888 2824 29952
rect 2888 29888 2896 29952
rect 1715 29204 1781 29205
rect 1715 29140 1716 29204
rect 1780 29140 1781 29204
rect 1715 29139 1781 29140
rect 2575 28864 2896 29888
rect 4207 31584 4527 32608
rect 4207 31520 4215 31584
rect 4279 31520 4295 31584
rect 4359 31520 4375 31584
rect 4439 31520 4455 31584
rect 4519 31520 4527 31584
rect 4207 30496 4527 31520
rect 4207 30432 4215 30496
rect 4279 30432 4295 30496
rect 4359 30432 4375 30496
rect 4439 30432 4455 30496
rect 4519 30432 4527 30496
rect 4207 29408 4527 30432
rect 4207 29344 4215 29408
rect 4279 29344 4295 29408
rect 4359 29344 4375 29408
rect 4439 29344 4455 29408
rect 4519 29344 4527 29408
rect 3003 28932 3069 28933
rect 3003 28868 3004 28932
rect 3068 28868 3069 28932
rect 3003 28867 3069 28868
rect 2575 28800 2584 28864
rect 2648 28800 2664 28864
rect 2728 28800 2744 28864
rect 2808 28800 2824 28864
rect 2888 28800 2896 28864
rect 2575 27776 2896 28800
rect 2575 27712 2584 27776
rect 2648 27712 2664 27776
rect 2728 27712 2744 27776
rect 2808 27712 2824 27776
rect 2888 27712 2896 27776
rect 2575 26688 2896 27712
rect 3006 26757 3066 28867
rect 4207 28320 4527 29344
rect 4207 28256 4215 28320
rect 4279 28256 4295 28320
rect 4359 28256 4375 28320
rect 4439 28256 4455 28320
rect 4519 28256 4527 28320
rect 4207 27232 4527 28256
rect 4207 27168 4215 27232
rect 4279 27168 4295 27232
rect 4359 27168 4375 27232
rect 4439 27168 4455 27232
rect 4519 27168 4527 27232
rect 3003 26756 3069 26757
rect 3003 26692 3004 26756
rect 3068 26692 3069 26756
rect 3003 26691 3069 26692
rect 2575 26624 2584 26688
rect 2648 26624 2664 26688
rect 2728 26624 2744 26688
rect 2808 26624 2824 26688
rect 2888 26624 2896 26688
rect 2575 25600 2896 26624
rect 2575 25536 2584 25600
rect 2648 25536 2664 25600
rect 2728 25536 2744 25600
rect 2808 25536 2824 25600
rect 2888 25536 2896 25600
rect 2575 24512 2896 25536
rect 2575 24448 2584 24512
rect 2648 24448 2664 24512
rect 2728 24448 2744 24512
rect 2808 24448 2824 24512
rect 2888 24448 2896 24512
rect 2575 23424 2896 24448
rect 2575 23360 2584 23424
rect 2648 23360 2664 23424
rect 2728 23360 2744 23424
rect 2808 23360 2824 23424
rect 2888 23360 2896 23424
rect 2575 22336 2896 23360
rect 2575 22272 2584 22336
rect 2648 22272 2664 22336
rect 2728 22272 2744 22336
rect 2808 22272 2824 22336
rect 2888 22272 2896 22336
rect 2575 21248 2896 22272
rect 2575 21184 2584 21248
rect 2648 21184 2664 21248
rect 2728 21184 2744 21248
rect 2808 21184 2824 21248
rect 2888 21184 2896 21248
rect 2575 20160 2896 21184
rect 2575 20096 2584 20160
rect 2648 20096 2664 20160
rect 2728 20096 2744 20160
rect 2808 20096 2824 20160
rect 2888 20096 2896 20160
rect 2575 19072 2896 20096
rect 2575 19008 2584 19072
rect 2648 19008 2664 19072
rect 2728 19008 2744 19072
rect 2808 19008 2824 19072
rect 2888 19008 2896 19072
rect 2575 17984 2896 19008
rect 2575 17920 2584 17984
rect 2648 17920 2664 17984
rect 2728 17920 2744 17984
rect 2808 17920 2824 17984
rect 2888 17920 2896 17984
rect 2575 16896 2896 17920
rect 2575 16832 2584 16896
rect 2648 16832 2664 16896
rect 2728 16832 2744 16896
rect 2808 16832 2824 16896
rect 2888 16832 2896 16896
rect 2575 15808 2896 16832
rect 2575 15744 2584 15808
rect 2648 15744 2664 15808
rect 2728 15744 2744 15808
rect 2808 15744 2824 15808
rect 2888 15744 2896 15808
rect 2575 14720 2896 15744
rect 2575 14656 2584 14720
rect 2648 14656 2664 14720
rect 2728 14656 2744 14720
rect 2808 14656 2824 14720
rect 2888 14656 2896 14720
rect 2575 13632 2896 14656
rect 2575 13568 2584 13632
rect 2648 13568 2664 13632
rect 2728 13568 2744 13632
rect 2808 13568 2824 13632
rect 2888 13568 2896 13632
rect 2575 12544 2896 13568
rect 2575 12480 2584 12544
rect 2648 12480 2664 12544
rect 2728 12480 2744 12544
rect 2808 12480 2824 12544
rect 2888 12480 2896 12544
rect 2575 11456 2896 12480
rect 2575 11392 2584 11456
rect 2648 11392 2664 11456
rect 2728 11392 2744 11456
rect 2808 11392 2824 11456
rect 2888 11392 2896 11456
rect 2575 10368 2896 11392
rect 2575 10304 2584 10368
rect 2648 10304 2664 10368
rect 2728 10304 2744 10368
rect 2808 10304 2824 10368
rect 2888 10304 2896 10368
rect 2575 9280 2896 10304
rect 2575 9216 2584 9280
rect 2648 9216 2664 9280
rect 2728 9216 2744 9280
rect 2808 9216 2824 9280
rect 2888 9216 2896 9280
rect 2575 8192 2896 9216
rect 2575 8128 2584 8192
rect 2648 8128 2664 8192
rect 2728 8128 2744 8192
rect 2808 8128 2824 8192
rect 2888 8128 2896 8192
rect 2575 7104 2896 8128
rect 2575 7040 2584 7104
rect 2648 7040 2664 7104
rect 2728 7040 2744 7104
rect 2808 7040 2824 7104
rect 2888 7040 2896 7104
rect 2575 6016 2896 7040
rect 2575 5952 2584 6016
rect 2648 5952 2664 6016
rect 2728 5952 2744 6016
rect 2808 5952 2824 6016
rect 2888 5952 2896 6016
rect 2575 4928 2896 5952
rect 2575 4864 2584 4928
rect 2648 4864 2664 4928
rect 2728 4864 2744 4928
rect 2808 4864 2824 4928
rect 2888 4864 2896 4928
rect 2575 3840 2896 4864
rect 2575 3776 2584 3840
rect 2648 3776 2664 3840
rect 2728 3776 2744 3840
rect 2808 3776 2824 3840
rect 2888 3776 2896 3840
rect 2575 2752 2896 3776
rect 2575 2688 2584 2752
rect 2648 2688 2664 2752
rect 2728 2688 2744 2752
rect 2808 2688 2824 2752
rect 2888 2688 2896 2752
rect 2575 2128 2896 2688
rect 4207 26144 4527 27168
rect 4207 26080 4215 26144
rect 4279 26080 4295 26144
rect 4359 26080 4375 26144
rect 4439 26080 4455 26144
rect 4519 26080 4527 26144
rect 4207 25056 4527 26080
rect 4207 24992 4215 25056
rect 4279 24992 4295 25056
rect 4359 24992 4375 25056
rect 4439 24992 4455 25056
rect 4519 24992 4527 25056
rect 4207 23968 4527 24992
rect 4207 23904 4215 23968
rect 4279 23904 4295 23968
rect 4359 23904 4375 23968
rect 4439 23904 4455 23968
rect 4519 23904 4527 23968
rect 4207 22880 4527 23904
rect 4207 22816 4215 22880
rect 4279 22816 4295 22880
rect 4359 22816 4375 22880
rect 4439 22816 4455 22880
rect 4519 22816 4527 22880
rect 4207 21792 4527 22816
rect 4207 21728 4215 21792
rect 4279 21728 4295 21792
rect 4359 21728 4375 21792
rect 4439 21728 4455 21792
rect 4519 21728 4527 21792
rect 4207 20704 4527 21728
rect 4207 20640 4215 20704
rect 4279 20640 4295 20704
rect 4359 20640 4375 20704
rect 4439 20640 4455 20704
rect 4519 20640 4527 20704
rect 4207 19616 4527 20640
rect 4207 19552 4215 19616
rect 4279 19552 4295 19616
rect 4359 19552 4375 19616
rect 4439 19552 4455 19616
rect 4519 19552 4527 19616
rect 4207 18528 4527 19552
rect 4207 18464 4215 18528
rect 4279 18464 4295 18528
rect 4359 18464 4375 18528
rect 4439 18464 4455 18528
rect 4519 18464 4527 18528
rect 4207 17440 4527 18464
rect 4207 17376 4215 17440
rect 4279 17376 4295 17440
rect 4359 17376 4375 17440
rect 4439 17376 4455 17440
rect 4519 17376 4527 17440
rect 4207 16352 4527 17376
rect 4207 16288 4215 16352
rect 4279 16288 4295 16352
rect 4359 16288 4375 16352
rect 4439 16288 4455 16352
rect 4519 16288 4527 16352
rect 4207 15264 4527 16288
rect 4207 15200 4215 15264
rect 4279 15200 4295 15264
rect 4359 15200 4375 15264
rect 4439 15200 4455 15264
rect 4519 15200 4527 15264
rect 4207 14176 4527 15200
rect 4207 14112 4215 14176
rect 4279 14112 4295 14176
rect 4359 14112 4375 14176
rect 4439 14112 4455 14176
rect 4519 14112 4527 14176
rect 4207 13088 4527 14112
rect 4207 13024 4215 13088
rect 4279 13024 4295 13088
rect 4359 13024 4375 13088
rect 4439 13024 4455 13088
rect 4519 13024 4527 13088
rect 4207 12000 4527 13024
rect 4207 11936 4215 12000
rect 4279 11936 4295 12000
rect 4359 11936 4375 12000
rect 4439 11936 4455 12000
rect 4519 11936 4527 12000
rect 4207 10912 4527 11936
rect 4207 10848 4215 10912
rect 4279 10848 4295 10912
rect 4359 10848 4375 10912
rect 4439 10848 4455 10912
rect 4519 10848 4527 10912
rect 4207 9824 4527 10848
rect 4207 9760 4215 9824
rect 4279 9760 4295 9824
rect 4359 9760 4375 9824
rect 4439 9760 4455 9824
rect 4519 9760 4527 9824
rect 4207 8736 4527 9760
rect 4207 8672 4215 8736
rect 4279 8672 4295 8736
rect 4359 8672 4375 8736
rect 4439 8672 4455 8736
rect 4519 8672 4527 8736
rect 4207 7648 4527 8672
rect 4207 7584 4215 7648
rect 4279 7584 4295 7648
rect 4359 7584 4375 7648
rect 4439 7584 4455 7648
rect 4519 7584 4527 7648
rect 4207 6560 4527 7584
rect 4207 6496 4215 6560
rect 4279 6496 4295 6560
rect 4359 6496 4375 6560
rect 4439 6496 4455 6560
rect 4519 6496 4527 6560
rect 4207 5472 4527 6496
rect 4207 5408 4215 5472
rect 4279 5408 4295 5472
rect 4359 5408 4375 5472
rect 4439 5408 4455 5472
rect 4519 5408 4527 5472
rect 4207 4384 4527 5408
rect 4207 4320 4215 4384
rect 4279 4320 4295 4384
rect 4359 4320 4375 4384
rect 4439 4320 4455 4384
rect 4519 4320 4527 4384
rect 4207 3296 4527 4320
rect 4207 3232 4215 3296
rect 4279 3232 4295 3296
rect 4359 3232 4375 3296
rect 4439 3232 4455 3296
rect 4519 3232 4527 3296
rect 4207 2208 4527 3232
rect 4207 2144 4215 2208
rect 4279 2144 4295 2208
rect 4359 2144 4375 2208
rect 4439 2144 4455 2208
rect 4519 2144 4527 2208
rect 4207 2128 4527 2144
rect 5839 38656 6159 39680
rect 5839 38592 5847 38656
rect 5911 38592 5927 38656
rect 5991 38592 6007 38656
rect 6071 38592 6087 38656
rect 6151 38592 6159 38656
rect 5839 37568 6159 38592
rect 5839 37504 5847 37568
rect 5911 37504 5927 37568
rect 5991 37504 6007 37568
rect 6071 37504 6087 37568
rect 6151 37504 6159 37568
rect 5839 36480 6159 37504
rect 5839 36416 5847 36480
rect 5911 36416 5927 36480
rect 5991 36416 6007 36480
rect 6071 36416 6087 36480
rect 6151 36416 6159 36480
rect 5839 35392 6159 36416
rect 5839 35328 5847 35392
rect 5911 35328 5927 35392
rect 5991 35328 6007 35392
rect 6071 35328 6087 35392
rect 6151 35328 6159 35392
rect 5839 34304 6159 35328
rect 5839 34240 5847 34304
rect 5911 34240 5927 34304
rect 5991 34240 6007 34304
rect 6071 34240 6087 34304
rect 6151 34240 6159 34304
rect 5839 33216 6159 34240
rect 5839 33152 5847 33216
rect 5911 33152 5927 33216
rect 5991 33152 6007 33216
rect 6071 33152 6087 33216
rect 6151 33152 6159 33216
rect 5839 32128 6159 33152
rect 5839 32064 5847 32128
rect 5911 32064 5927 32128
rect 5991 32064 6007 32128
rect 6071 32064 6087 32128
rect 6151 32064 6159 32128
rect 5839 31040 6159 32064
rect 5839 30976 5847 31040
rect 5911 30976 5927 31040
rect 5991 30976 6007 31040
rect 6071 30976 6087 31040
rect 6151 30976 6159 31040
rect 5839 29952 6159 30976
rect 5839 29888 5847 29952
rect 5911 29888 5927 29952
rect 5991 29888 6007 29952
rect 6071 29888 6087 29952
rect 6151 29888 6159 29952
rect 5839 28864 6159 29888
rect 5839 28800 5847 28864
rect 5911 28800 5927 28864
rect 5991 28800 6007 28864
rect 6071 28800 6087 28864
rect 6151 28800 6159 28864
rect 5839 27776 6159 28800
rect 5839 27712 5847 27776
rect 5911 27712 5927 27776
rect 5991 27712 6007 27776
rect 6071 27712 6087 27776
rect 6151 27712 6159 27776
rect 5839 26688 6159 27712
rect 5839 26624 5847 26688
rect 5911 26624 5927 26688
rect 5991 26624 6007 26688
rect 6071 26624 6087 26688
rect 6151 26624 6159 26688
rect 5839 25600 6159 26624
rect 5839 25536 5847 25600
rect 5911 25536 5927 25600
rect 5991 25536 6007 25600
rect 6071 25536 6087 25600
rect 6151 25536 6159 25600
rect 5839 24512 6159 25536
rect 5839 24448 5847 24512
rect 5911 24448 5927 24512
rect 5991 24448 6007 24512
rect 6071 24448 6087 24512
rect 6151 24448 6159 24512
rect 5839 23424 6159 24448
rect 5839 23360 5847 23424
rect 5911 23360 5927 23424
rect 5991 23360 6007 23424
rect 6071 23360 6087 23424
rect 6151 23360 6159 23424
rect 5839 22336 6159 23360
rect 5839 22272 5847 22336
rect 5911 22272 5927 22336
rect 5991 22272 6007 22336
rect 6071 22272 6087 22336
rect 6151 22272 6159 22336
rect 5839 21248 6159 22272
rect 5839 21184 5847 21248
rect 5911 21184 5927 21248
rect 5991 21184 6007 21248
rect 6071 21184 6087 21248
rect 6151 21184 6159 21248
rect 5839 20160 6159 21184
rect 5839 20096 5847 20160
rect 5911 20096 5927 20160
rect 5991 20096 6007 20160
rect 6071 20096 6087 20160
rect 6151 20096 6159 20160
rect 5839 19072 6159 20096
rect 5839 19008 5847 19072
rect 5911 19008 5927 19072
rect 5991 19008 6007 19072
rect 6071 19008 6087 19072
rect 6151 19008 6159 19072
rect 5839 17984 6159 19008
rect 5839 17920 5847 17984
rect 5911 17920 5927 17984
rect 5991 17920 6007 17984
rect 6071 17920 6087 17984
rect 6151 17920 6159 17984
rect 5839 16896 6159 17920
rect 5839 16832 5847 16896
rect 5911 16832 5927 16896
rect 5991 16832 6007 16896
rect 6071 16832 6087 16896
rect 6151 16832 6159 16896
rect 5839 15808 6159 16832
rect 5839 15744 5847 15808
rect 5911 15744 5927 15808
rect 5991 15744 6007 15808
rect 6071 15744 6087 15808
rect 6151 15744 6159 15808
rect 5839 14720 6159 15744
rect 5839 14656 5847 14720
rect 5911 14656 5927 14720
rect 5991 14656 6007 14720
rect 6071 14656 6087 14720
rect 6151 14656 6159 14720
rect 5839 13632 6159 14656
rect 5839 13568 5847 13632
rect 5911 13568 5927 13632
rect 5991 13568 6007 13632
rect 6071 13568 6087 13632
rect 6151 13568 6159 13632
rect 5839 12544 6159 13568
rect 5839 12480 5847 12544
rect 5911 12480 5927 12544
rect 5991 12480 6007 12544
rect 6071 12480 6087 12544
rect 6151 12480 6159 12544
rect 5839 11456 6159 12480
rect 5839 11392 5847 11456
rect 5911 11392 5927 11456
rect 5991 11392 6007 11456
rect 6071 11392 6087 11456
rect 6151 11392 6159 11456
rect 5839 10368 6159 11392
rect 5839 10304 5847 10368
rect 5911 10304 5927 10368
rect 5991 10304 6007 10368
rect 6071 10304 6087 10368
rect 6151 10304 6159 10368
rect 5839 9280 6159 10304
rect 5839 9216 5847 9280
rect 5911 9216 5927 9280
rect 5991 9216 6007 9280
rect 6071 9216 6087 9280
rect 6151 9216 6159 9280
rect 5839 8192 6159 9216
rect 5839 8128 5847 8192
rect 5911 8128 5927 8192
rect 5991 8128 6007 8192
rect 6071 8128 6087 8192
rect 6151 8128 6159 8192
rect 5839 7104 6159 8128
rect 5839 7040 5847 7104
rect 5911 7040 5927 7104
rect 5991 7040 6007 7104
rect 6071 7040 6087 7104
rect 6151 7040 6159 7104
rect 5839 6016 6159 7040
rect 5839 5952 5847 6016
rect 5911 5952 5927 6016
rect 5991 5952 6007 6016
rect 6071 5952 6087 6016
rect 6151 5952 6159 6016
rect 5839 4928 6159 5952
rect 5839 4864 5847 4928
rect 5911 4864 5927 4928
rect 5991 4864 6007 4928
rect 6071 4864 6087 4928
rect 6151 4864 6159 4928
rect 5839 3840 6159 4864
rect 5839 3776 5847 3840
rect 5911 3776 5927 3840
rect 5991 3776 6007 3840
rect 6071 3776 6087 3840
rect 6151 3776 6159 3840
rect 5839 2752 6159 3776
rect 5839 2688 5847 2752
rect 5911 2688 5927 2752
rect 5991 2688 6007 2752
rect 6071 2688 6087 2752
rect 6151 2688 6159 2752
rect 5839 2128 6159 2688
rect 7471 40288 7791 41312
rect 7471 40224 7479 40288
rect 7543 40224 7559 40288
rect 7623 40224 7639 40288
rect 7703 40224 7719 40288
rect 7783 40224 7791 40288
rect 7471 39200 7791 40224
rect 7471 39136 7479 39200
rect 7543 39136 7559 39200
rect 7623 39136 7639 39200
rect 7703 39136 7719 39200
rect 7783 39136 7791 39200
rect 7471 38112 7791 39136
rect 7471 38048 7479 38112
rect 7543 38048 7559 38112
rect 7623 38048 7639 38112
rect 7703 38048 7719 38112
rect 7783 38048 7791 38112
rect 7471 37024 7791 38048
rect 7471 36960 7479 37024
rect 7543 36960 7559 37024
rect 7623 36960 7639 37024
rect 7703 36960 7719 37024
rect 7783 36960 7791 37024
rect 7471 35936 7791 36960
rect 7471 35872 7479 35936
rect 7543 35872 7559 35936
rect 7623 35872 7639 35936
rect 7703 35872 7719 35936
rect 7783 35872 7791 35936
rect 7471 34848 7791 35872
rect 7471 34784 7479 34848
rect 7543 34784 7559 34848
rect 7623 34784 7639 34848
rect 7703 34784 7719 34848
rect 7783 34784 7791 34848
rect 7471 33760 7791 34784
rect 7471 33696 7479 33760
rect 7543 33696 7559 33760
rect 7623 33696 7639 33760
rect 7703 33696 7719 33760
rect 7783 33696 7791 33760
rect 7471 32672 7791 33696
rect 7471 32608 7479 32672
rect 7543 32608 7559 32672
rect 7623 32608 7639 32672
rect 7703 32608 7719 32672
rect 7783 32608 7791 32672
rect 7471 31584 7791 32608
rect 7471 31520 7479 31584
rect 7543 31520 7559 31584
rect 7623 31520 7639 31584
rect 7703 31520 7719 31584
rect 7783 31520 7791 31584
rect 7471 30496 7791 31520
rect 7471 30432 7479 30496
rect 7543 30432 7559 30496
rect 7623 30432 7639 30496
rect 7703 30432 7719 30496
rect 7783 30432 7791 30496
rect 7471 29408 7791 30432
rect 7471 29344 7479 29408
rect 7543 29344 7559 29408
rect 7623 29344 7639 29408
rect 7703 29344 7719 29408
rect 7783 29344 7791 29408
rect 7471 28320 7791 29344
rect 7471 28256 7479 28320
rect 7543 28256 7559 28320
rect 7623 28256 7639 28320
rect 7703 28256 7719 28320
rect 7783 28256 7791 28320
rect 7471 27232 7791 28256
rect 7471 27168 7479 27232
rect 7543 27168 7559 27232
rect 7623 27168 7639 27232
rect 7703 27168 7719 27232
rect 7783 27168 7791 27232
rect 7471 26144 7791 27168
rect 7471 26080 7479 26144
rect 7543 26080 7559 26144
rect 7623 26080 7639 26144
rect 7703 26080 7719 26144
rect 7783 26080 7791 26144
rect 7471 25056 7791 26080
rect 7471 24992 7479 25056
rect 7543 24992 7559 25056
rect 7623 24992 7639 25056
rect 7703 24992 7719 25056
rect 7783 24992 7791 25056
rect 7471 23968 7791 24992
rect 7471 23904 7479 23968
rect 7543 23904 7559 23968
rect 7623 23904 7639 23968
rect 7703 23904 7719 23968
rect 7783 23904 7791 23968
rect 7471 22880 7791 23904
rect 7471 22816 7479 22880
rect 7543 22816 7559 22880
rect 7623 22816 7639 22880
rect 7703 22816 7719 22880
rect 7783 22816 7791 22880
rect 7471 21792 7791 22816
rect 7471 21728 7479 21792
rect 7543 21728 7559 21792
rect 7623 21728 7639 21792
rect 7703 21728 7719 21792
rect 7783 21728 7791 21792
rect 7471 20704 7791 21728
rect 7471 20640 7479 20704
rect 7543 20640 7559 20704
rect 7623 20640 7639 20704
rect 7703 20640 7719 20704
rect 7783 20640 7791 20704
rect 7471 19616 7791 20640
rect 7471 19552 7479 19616
rect 7543 19552 7559 19616
rect 7623 19552 7639 19616
rect 7703 19552 7719 19616
rect 7783 19552 7791 19616
rect 7471 18528 7791 19552
rect 7471 18464 7479 18528
rect 7543 18464 7559 18528
rect 7623 18464 7639 18528
rect 7703 18464 7719 18528
rect 7783 18464 7791 18528
rect 7471 17440 7791 18464
rect 7471 17376 7479 17440
rect 7543 17376 7559 17440
rect 7623 17376 7639 17440
rect 7703 17376 7719 17440
rect 7783 17376 7791 17440
rect 7471 16352 7791 17376
rect 7471 16288 7479 16352
rect 7543 16288 7559 16352
rect 7623 16288 7639 16352
rect 7703 16288 7719 16352
rect 7783 16288 7791 16352
rect 7471 15264 7791 16288
rect 7471 15200 7479 15264
rect 7543 15200 7559 15264
rect 7623 15200 7639 15264
rect 7703 15200 7719 15264
rect 7783 15200 7791 15264
rect 7471 14176 7791 15200
rect 7471 14112 7479 14176
rect 7543 14112 7559 14176
rect 7623 14112 7639 14176
rect 7703 14112 7719 14176
rect 7783 14112 7791 14176
rect 7471 13088 7791 14112
rect 7471 13024 7479 13088
rect 7543 13024 7559 13088
rect 7623 13024 7639 13088
rect 7703 13024 7719 13088
rect 7783 13024 7791 13088
rect 7471 12000 7791 13024
rect 7471 11936 7479 12000
rect 7543 11936 7559 12000
rect 7623 11936 7639 12000
rect 7703 11936 7719 12000
rect 7783 11936 7791 12000
rect 7471 10912 7791 11936
rect 7471 10848 7479 10912
rect 7543 10848 7559 10912
rect 7623 10848 7639 10912
rect 7703 10848 7719 10912
rect 7783 10848 7791 10912
rect 7471 9824 7791 10848
rect 7471 9760 7479 9824
rect 7543 9760 7559 9824
rect 7623 9760 7639 9824
rect 7703 9760 7719 9824
rect 7783 9760 7791 9824
rect 7471 8736 7791 9760
rect 7471 8672 7479 8736
rect 7543 8672 7559 8736
rect 7623 8672 7639 8736
rect 7703 8672 7719 8736
rect 7783 8672 7791 8736
rect 7471 7648 7791 8672
rect 7471 7584 7479 7648
rect 7543 7584 7559 7648
rect 7623 7584 7639 7648
rect 7703 7584 7719 7648
rect 7783 7584 7791 7648
rect 7471 6560 7791 7584
rect 7471 6496 7479 6560
rect 7543 6496 7559 6560
rect 7623 6496 7639 6560
rect 7703 6496 7719 6560
rect 7783 6496 7791 6560
rect 7471 5472 7791 6496
rect 7471 5408 7479 5472
rect 7543 5408 7559 5472
rect 7623 5408 7639 5472
rect 7703 5408 7719 5472
rect 7783 5408 7791 5472
rect 7471 4384 7791 5408
rect 7471 4320 7479 4384
rect 7543 4320 7559 4384
rect 7623 4320 7639 4384
rect 7703 4320 7719 4384
rect 7783 4320 7791 4384
rect 7471 3296 7791 4320
rect 7471 3232 7479 3296
rect 7543 3232 7559 3296
rect 7623 3232 7639 3296
rect 7703 3232 7719 3296
rect 7783 3232 7791 3296
rect 7471 2208 7791 3232
rect 7471 2144 7479 2208
rect 7543 2144 7559 2208
rect 7623 2144 7639 2208
rect 7703 2144 7719 2208
rect 7783 2144 7791 2208
rect 7471 2128 7791 2144
rect 9103 77824 9423 77840
rect 9103 77760 9111 77824
rect 9175 77760 9191 77824
rect 9255 77760 9271 77824
rect 9335 77760 9351 77824
rect 9415 77760 9423 77824
rect 9103 76736 9423 77760
rect 9103 76672 9111 76736
rect 9175 76672 9191 76736
rect 9255 76672 9271 76736
rect 9335 76672 9351 76736
rect 9415 76672 9423 76736
rect 9103 75648 9423 76672
rect 9103 75584 9111 75648
rect 9175 75584 9191 75648
rect 9255 75584 9271 75648
rect 9335 75584 9351 75648
rect 9415 75584 9423 75648
rect 9103 74560 9423 75584
rect 9103 74496 9111 74560
rect 9175 74496 9191 74560
rect 9255 74496 9271 74560
rect 9335 74496 9351 74560
rect 9415 74496 9423 74560
rect 9103 73472 9423 74496
rect 9103 73408 9111 73472
rect 9175 73408 9191 73472
rect 9255 73408 9271 73472
rect 9335 73408 9351 73472
rect 9415 73408 9423 73472
rect 9103 72384 9423 73408
rect 9103 72320 9111 72384
rect 9175 72320 9191 72384
rect 9255 72320 9271 72384
rect 9335 72320 9351 72384
rect 9415 72320 9423 72384
rect 9103 71296 9423 72320
rect 9103 71232 9111 71296
rect 9175 71232 9191 71296
rect 9255 71232 9271 71296
rect 9335 71232 9351 71296
rect 9415 71232 9423 71296
rect 9103 70208 9423 71232
rect 9103 70144 9111 70208
rect 9175 70144 9191 70208
rect 9255 70144 9271 70208
rect 9335 70144 9351 70208
rect 9415 70144 9423 70208
rect 9103 69120 9423 70144
rect 9103 69056 9111 69120
rect 9175 69056 9191 69120
rect 9255 69056 9271 69120
rect 9335 69056 9351 69120
rect 9415 69056 9423 69120
rect 9103 68032 9423 69056
rect 9103 67968 9111 68032
rect 9175 67968 9191 68032
rect 9255 67968 9271 68032
rect 9335 67968 9351 68032
rect 9415 67968 9423 68032
rect 9103 66944 9423 67968
rect 9103 66880 9111 66944
rect 9175 66880 9191 66944
rect 9255 66880 9271 66944
rect 9335 66880 9351 66944
rect 9415 66880 9423 66944
rect 9103 65856 9423 66880
rect 9103 65792 9111 65856
rect 9175 65792 9191 65856
rect 9255 65792 9271 65856
rect 9335 65792 9351 65856
rect 9415 65792 9423 65856
rect 9103 64768 9423 65792
rect 9103 64704 9111 64768
rect 9175 64704 9191 64768
rect 9255 64704 9271 64768
rect 9335 64704 9351 64768
rect 9415 64704 9423 64768
rect 9103 63680 9423 64704
rect 9103 63616 9111 63680
rect 9175 63616 9191 63680
rect 9255 63616 9271 63680
rect 9335 63616 9351 63680
rect 9415 63616 9423 63680
rect 9103 62592 9423 63616
rect 9103 62528 9111 62592
rect 9175 62528 9191 62592
rect 9255 62528 9271 62592
rect 9335 62528 9351 62592
rect 9415 62528 9423 62592
rect 9103 61504 9423 62528
rect 9103 61440 9111 61504
rect 9175 61440 9191 61504
rect 9255 61440 9271 61504
rect 9335 61440 9351 61504
rect 9415 61440 9423 61504
rect 9103 60416 9423 61440
rect 9103 60352 9111 60416
rect 9175 60352 9191 60416
rect 9255 60352 9271 60416
rect 9335 60352 9351 60416
rect 9415 60352 9423 60416
rect 9103 59328 9423 60352
rect 9103 59264 9111 59328
rect 9175 59264 9191 59328
rect 9255 59264 9271 59328
rect 9335 59264 9351 59328
rect 9415 59264 9423 59328
rect 9103 58240 9423 59264
rect 9103 58176 9111 58240
rect 9175 58176 9191 58240
rect 9255 58176 9271 58240
rect 9335 58176 9351 58240
rect 9415 58176 9423 58240
rect 9103 57152 9423 58176
rect 9103 57088 9111 57152
rect 9175 57088 9191 57152
rect 9255 57088 9271 57152
rect 9335 57088 9351 57152
rect 9415 57088 9423 57152
rect 9103 56064 9423 57088
rect 9103 56000 9111 56064
rect 9175 56000 9191 56064
rect 9255 56000 9271 56064
rect 9335 56000 9351 56064
rect 9415 56000 9423 56064
rect 9103 54976 9423 56000
rect 9103 54912 9111 54976
rect 9175 54912 9191 54976
rect 9255 54912 9271 54976
rect 9335 54912 9351 54976
rect 9415 54912 9423 54976
rect 9103 53888 9423 54912
rect 9103 53824 9111 53888
rect 9175 53824 9191 53888
rect 9255 53824 9271 53888
rect 9335 53824 9351 53888
rect 9415 53824 9423 53888
rect 9103 52800 9423 53824
rect 9103 52736 9111 52800
rect 9175 52736 9191 52800
rect 9255 52736 9271 52800
rect 9335 52736 9351 52800
rect 9415 52736 9423 52800
rect 9103 51712 9423 52736
rect 9103 51648 9111 51712
rect 9175 51648 9191 51712
rect 9255 51648 9271 51712
rect 9335 51648 9351 51712
rect 9415 51648 9423 51712
rect 9103 50624 9423 51648
rect 9103 50560 9111 50624
rect 9175 50560 9191 50624
rect 9255 50560 9271 50624
rect 9335 50560 9351 50624
rect 9415 50560 9423 50624
rect 9103 49536 9423 50560
rect 9103 49472 9111 49536
rect 9175 49472 9191 49536
rect 9255 49472 9271 49536
rect 9335 49472 9351 49536
rect 9415 49472 9423 49536
rect 9103 48448 9423 49472
rect 9103 48384 9111 48448
rect 9175 48384 9191 48448
rect 9255 48384 9271 48448
rect 9335 48384 9351 48448
rect 9415 48384 9423 48448
rect 9103 47360 9423 48384
rect 9103 47296 9111 47360
rect 9175 47296 9191 47360
rect 9255 47296 9271 47360
rect 9335 47296 9351 47360
rect 9415 47296 9423 47360
rect 9103 46272 9423 47296
rect 9103 46208 9111 46272
rect 9175 46208 9191 46272
rect 9255 46208 9271 46272
rect 9335 46208 9351 46272
rect 9415 46208 9423 46272
rect 9103 45184 9423 46208
rect 9103 45120 9111 45184
rect 9175 45120 9191 45184
rect 9255 45120 9271 45184
rect 9335 45120 9351 45184
rect 9415 45120 9423 45184
rect 9103 44096 9423 45120
rect 9103 44032 9111 44096
rect 9175 44032 9191 44096
rect 9255 44032 9271 44096
rect 9335 44032 9351 44096
rect 9415 44032 9423 44096
rect 9103 43008 9423 44032
rect 9103 42944 9111 43008
rect 9175 42944 9191 43008
rect 9255 42944 9271 43008
rect 9335 42944 9351 43008
rect 9415 42944 9423 43008
rect 9103 41920 9423 42944
rect 9103 41856 9111 41920
rect 9175 41856 9191 41920
rect 9255 41856 9271 41920
rect 9335 41856 9351 41920
rect 9415 41856 9423 41920
rect 9103 40832 9423 41856
rect 9103 40768 9111 40832
rect 9175 40768 9191 40832
rect 9255 40768 9271 40832
rect 9335 40768 9351 40832
rect 9415 40768 9423 40832
rect 9103 39744 9423 40768
rect 9103 39680 9111 39744
rect 9175 39680 9191 39744
rect 9255 39680 9271 39744
rect 9335 39680 9351 39744
rect 9415 39680 9423 39744
rect 9103 38656 9423 39680
rect 9103 38592 9111 38656
rect 9175 38592 9191 38656
rect 9255 38592 9271 38656
rect 9335 38592 9351 38656
rect 9415 38592 9423 38656
rect 9103 37568 9423 38592
rect 9103 37504 9111 37568
rect 9175 37504 9191 37568
rect 9255 37504 9271 37568
rect 9335 37504 9351 37568
rect 9415 37504 9423 37568
rect 9103 36480 9423 37504
rect 9103 36416 9111 36480
rect 9175 36416 9191 36480
rect 9255 36416 9271 36480
rect 9335 36416 9351 36480
rect 9415 36416 9423 36480
rect 9103 35392 9423 36416
rect 9103 35328 9111 35392
rect 9175 35328 9191 35392
rect 9255 35328 9271 35392
rect 9335 35328 9351 35392
rect 9415 35328 9423 35392
rect 9103 34304 9423 35328
rect 9103 34240 9111 34304
rect 9175 34240 9191 34304
rect 9255 34240 9271 34304
rect 9335 34240 9351 34304
rect 9415 34240 9423 34304
rect 9103 33216 9423 34240
rect 9103 33152 9111 33216
rect 9175 33152 9191 33216
rect 9255 33152 9271 33216
rect 9335 33152 9351 33216
rect 9415 33152 9423 33216
rect 9103 32128 9423 33152
rect 9103 32064 9111 32128
rect 9175 32064 9191 32128
rect 9255 32064 9271 32128
rect 9335 32064 9351 32128
rect 9415 32064 9423 32128
rect 9103 31040 9423 32064
rect 9103 30976 9111 31040
rect 9175 30976 9191 31040
rect 9255 30976 9271 31040
rect 9335 30976 9351 31040
rect 9415 30976 9423 31040
rect 9103 29952 9423 30976
rect 9103 29888 9111 29952
rect 9175 29888 9191 29952
rect 9255 29888 9271 29952
rect 9335 29888 9351 29952
rect 9415 29888 9423 29952
rect 9103 28864 9423 29888
rect 9103 28800 9111 28864
rect 9175 28800 9191 28864
rect 9255 28800 9271 28864
rect 9335 28800 9351 28864
rect 9415 28800 9423 28864
rect 9103 27776 9423 28800
rect 9103 27712 9111 27776
rect 9175 27712 9191 27776
rect 9255 27712 9271 27776
rect 9335 27712 9351 27776
rect 9415 27712 9423 27776
rect 9103 26688 9423 27712
rect 9103 26624 9111 26688
rect 9175 26624 9191 26688
rect 9255 26624 9271 26688
rect 9335 26624 9351 26688
rect 9415 26624 9423 26688
rect 9103 25600 9423 26624
rect 9103 25536 9111 25600
rect 9175 25536 9191 25600
rect 9255 25536 9271 25600
rect 9335 25536 9351 25600
rect 9415 25536 9423 25600
rect 9103 24512 9423 25536
rect 9103 24448 9111 24512
rect 9175 24448 9191 24512
rect 9255 24448 9271 24512
rect 9335 24448 9351 24512
rect 9415 24448 9423 24512
rect 9103 23424 9423 24448
rect 9103 23360 9111 23424
rect 9175 23360 9191 23424
rect 9255 23360 9271 23424
rect 9335 23360 9351 23424
rect 9415 23360 9423 23424
rect 9103 22336 9423 23360
rect 9103 22272 9111 22336
rect 9175 22272 9191 22336
rect 9255 22272 9271 22336
rect 9335 22272 9351 22336
rect 9415 22272 9423 22336
rect 9103 21248 9423 22272
rect 9103 21184 9111 21248
rect 9175 21184 9191 21248
rect 9255 21184 9271 21248
rect 9335 21184 9351 21248
rect 9415 21184 9423 21248
rect 9103 20160 9423 21184
rect 9103 20096 9111 20160
rect 9175 20096 9191 20160
rect 9255 20096 9271 20160
rect 9335 20096 9351 20160
rect 9415 20096 9423 20160
rect 9103 19072 9423 20096
rect 9103 19008 9111 19072
rect 9175 19008 9191 19072
rect 9255 19008 9271 19072
rect 9335 19008 9351 19072
rect 9415 19008 9423 19072
rect 9103 17984 9423 19008
rect 9103 17920 9111 17984
rect 9175 17920 9191 17984
rect 9255 17920 9271 17984
rect 9335 17920 9351 17984
rect 9415 17920 9423 17984
rect 9103 16896 9423 17920
rect 9103 16832 9111 16896
rect 9175 16832 9191 16896
rect 9255 16832 9271 16896
rect 9335 16832 9351 16896
rect 9415 16832 9423 16896
rect 9103 15808 9423 16832
rect 9103 15744 9111 15808
rect 9175 15744 9191 15808
rect 9255 15744 9271 15808
rect 9335 15744 9351 15808
rect 9415 15744 9423 15808
rect 9103 14720 9423 15744
rect 9103 14656 9111 14720
rect 9175 14656 9191 14720
rect 9255 14656 9271 14720
rect 9335 14656 9351 14720
rect 9415 14656 9423 14720
rect 9103 13632 9423 14656
rect 9103 13568 9111 13632
rect 9175 13568 9191 13632
rect 9255 13568 9271 13632
rect 9335 13568 9351 13632
rect 9415 13568 9423 13632
rect 9103 12544 9423 13568
rect 9103 12480 9111 12544
rect 9175 12480 9191 12544
rect 9255 12480 9271 12544
rect 9335 12480 9351 12544
rect 9415 12480 9423 12544
rect 9103 11456 9423 12480
rect 9103 11392 9111 11456
rect 9175 11392 9191 11456
rect 9255 11392 9271 11456
rect 9335 11392 9351 11456
rect 9415 11392 9423 11456
rect 9103 10368 9423 11392
rect 9103 10304 9111 10368
rect 9175 10304 9191 10368
rect 9255 10304 9271 10368
rect 9335 10304 9351 10368
rect 9415 10304 9423 10368
rect 9103 9280 9423 10304
rect 9103 9216 9111 9280
rect 9175 9216 9191 9280
rect 9255 9216 9271 9280
rect 9335 9216 9351 9280
rect 9415 9216 9423 9280
rect 9103 8192 9423 9216
rect 9103 8128 9111 8192
rect 9175 8128 9191 8192
rect 9255 8128 9271 8192
rect 9335 8128 9351 8192
rect 9415 8128 9423 8192
rect 9103 7104 9423 8128
rect 9103 7040 9111 7104
rect 9175 7040 9191 7104
rect 9255 7040 9271 7104
rect 9335 7040 9351 7104
rect 9415 7040 9423 7104
rect 9103 6016 9423 7040
rect 9103 5952 9111 6016
rect 9175 5952 9191 6016
rect 9255 5952 9271 6016
rect 9335 5952 9351 6016
rect 9415 5952 9423 6016
rect 9103 4928 9423 5952
rect 9103 4864 9111 4928
rect 9175 4864 9191 4928
rect 9255 4864 9271 4928
rect 9335 4864 9351 4928
rect 9415 4864 9423 4928
rect 9103 3840 9423 4864
rect 9103 3776 9111 3840
rect 9175 3776 9191 3840
rect 9255 3776 9271 3840
rect 9335 3776 9351 3840
rect 9415 3776 9423 3840
rect 9103 2752 9423 3776
rect 9103 2688 9111 2752
rect 9175 2688 9191 2752
rect 9255 2688 9271 2752
rect 9335 2688 9351 2752
rect 9415 2688 9423 2752
rect 9103 2128 9423 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1635444444
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input135 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1635444444
transform -1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13
timestamp 1635444444
transform 1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1635444444
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_20
timestamp 1635444444
transform 1 0 2944 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1635444444
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1635444444
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1635444444
transform 1 0 2668 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1635444444
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1635444444
transform 1 0 3588 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1635444444
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1635444444
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1635444444
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_39
timestamp 1635444444
transform 1 0 4692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51
timestamp 1635444444
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp 1635444444
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1635444444
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1635444444
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1635444444
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1635444444
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1635444444
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1635444444
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1635444444
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1635444444
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 8556 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1635444444
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output199 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1635444444
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91
timestamp 1635444444
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1635444444
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_91
timestamp 1635444444
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_99
timestamp 1635444444
transform 1 0 10212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1635444444
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1635444444
transform 1 0 9844 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1635444444
transform -1 0 10856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1635444444
transform -1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1635444444
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1635444444
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _316_
timestamp 1635444444
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_14
timestamp 1635444444
transform 1 0 2392 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1635444444
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 3220 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1635444444
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1635444444
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1635444444
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1635444444
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1635444444
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1635444444
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1635444444
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1635444444
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1635444444
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1635444444
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1635444444
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1635444444
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1635444444
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1635444444
transform -1 0 10856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1635444444
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1635444444
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1635444444
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1635444444
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1635444444
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _220_
timestamp 1635444444
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _221_
timestamp 1635444444
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1635444444
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_34
timestamp 1635444444
transform 1 0 4232 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1635444444
transform 1 0 3956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_46
timestamp 1635444444
transform 1 0 5336 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1635444444
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1635444444
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1635444444
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1635444444
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1635444444
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1635444444
transform 1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_93
timestamp 1635444444
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1635444444
transform -1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7
timestamp 1635444444
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1635444444
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _306_
timestamp 1635444444
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1635444444
transform 1 0 2300 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1635444444
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1635444444
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _281_
timestamp 1635444444
transform -1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _305_
timestamp 1635444444
transform -1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1635444444
transform 1 0 4048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1635444444
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1635444444
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1635444444
transform 1 0 5152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1635444444
transform 1 0 6256 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1635444444
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1635444444
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1635444444
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1635444444
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1635444444
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1635444444
transform 1 0 10212 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1635444444
transform 1 0 9844 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1635444444
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_11
timestamp 1635444444
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1635444444
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1635444444
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1635444444
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 1635444444
transform -1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1635444444
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_23
timestamp 1635444444
transform 1 0 3220 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _219_
timestamp 1635444444
transform -1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_35
timestamp 1635444444
transform 1 0 4324 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1635444444
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1635444444
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1635444444
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1635444444
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1635444444
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1635444444
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1635444444
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1635444444
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1635444444
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1635444444
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1635444444
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1635444444
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1635444444
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1635444444
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1635444444
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1635444444
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _214_
timestamp 1635444444
transform -1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _283_
timestamp 1635444444
transform -1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _307_
timestamp 1635444444
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_14
timestamp 1635444444
transform 1 0 2392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1635444444
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1635444444
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _282_
timestamp 1635444444
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1635444444
transform 1 0 2760 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1635444444
transform 1 0 3220 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1635444444
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1635444444
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1635444444
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1635444444
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1635444444
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1635444444
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1635444444
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1635444444
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1635444444
transform 1 0 6256 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1635444444
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1635444444
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1635444444
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1635444444
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1635444444
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1635444444
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1635444444
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1635444444
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1635444444
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1635444444
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1635444444
transform 1 0 10396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1635444444
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1635444444
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1635444444
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1635444444
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1635444444
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1635444444
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_13
timestamp 1635444444
transform 1 0 2300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1635444444
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _308_
timestamp 1635444444
transform -1 0 3036 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1635444444
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1635444444
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1635444444
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1635444444
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1635444444
transform 1 0 5152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1635444444
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1635444444
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1635444444
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1635444444
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1635444444
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1635444444
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1635444444
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1635444444
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1635444444
transform -1 0 10856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1635444444
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1635444444
transform 1 0 1380 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_9_13
timestamp 1635444444
transform 1 0 2300 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_21
timestamp 1635444444
transform 1 0 3036 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _225_
timestamp 1635444444
transform -1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input98
timestamp 1635444444
transform 1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_28
timestamp 1635444444
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_40
timestamp 1635444444
transform 1 0 4784 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1635444444
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1635444444
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1635444444
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1635444444
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1635444444
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1635444444
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1635444444
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1635444444
transform 1 0 9844 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1635444444
transform -1 0 10856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1635444444
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1635444444
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_8  FILLER_10_13
timestamp 1635444444
transform 1 0 2300 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1635444444
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _217_
timestamp 1635444444
transform -1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1635444444
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1635444444
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1635444444
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1635444444
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1635444444
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1635444444
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1635444444
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1635444444
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1635444444
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_97
timestamp 1635444444
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1635444444
transform -1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_6
timestamp 1635444444
transform 1 0 1656 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1635444444
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1635444444
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_14
timestamp 1635444444
transform 1 0 2392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_18
timestamp 1635444444
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _284_
timestamp 1635444444
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1635444444
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1635444444
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1635444444
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1635444444
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1635444444
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1635444444
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_81
timestamp 1635444444
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 1635444444
transform 1 0 9108 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _294_
timestamp 1635444444
transform -1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_91
timestamp 1635444444
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1635444444
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1635444444
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1635444444
transform -1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1635444444
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_8
timestamp 1635444444
transform 1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1635444444
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _285_
timestamp 1635444444
transform -1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _310_
timestamp 1635444444
transform -1 0 1840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1635444444
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1635444444
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _286_
timestamp 1635444444
transform -1 0 3128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1635444444
transform 1 0 4048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1635444444
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1635444444
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1635444444
transform 1 0 5152 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1635444444
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1635444444
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1635444444
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1635444444
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1635444444
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1635444444
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_91
timestamp 1635444444
transform 1 0 9476 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1635444444
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1635444444
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1635444444
transform -1 0 10856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1635444444
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1635444444
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1635444444
transform 1 0 1380 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1635444444
transform 1 0 1380 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1635444444
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_22
timestamp 1635444444
transform 1 0 3128 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_13
timestamp 1635444444
transform 1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1635444444
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _087_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2668 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _309_
timestamp 1635444444
transform -1 0 3036 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_34
timestamp 1635444444
transform 1 0 4232 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1635444444
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1635444444
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1635444444
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1635444444
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1635444444
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1635444444
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1635444444
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1635444444
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1635444444
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1635444444
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1635444444
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1635444444
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1635444444
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1635444444
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1635444444
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1635444444
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_93
timestamp 1635444444
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_99
timestamp 1635444444
transform 1 0 10212 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1635444444
transform 1 0 10028 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1635444444
transform 1 0 9844 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1635444444
transform -1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1635444444
transform -1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1635444444
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1635444444
transform 1 0 1380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1635444444
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_20
timestamp 1635444444
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _287_
timestamp 1635444444
transform -1 0 2944 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1635444444
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1635444444
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1635444444
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1635444444
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1635444444
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1635444444
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1635444444
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1635444444
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1635444444
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1635444444
transform -1 0 10856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1635444444
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1635444444
transform 1 0 1380 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_16_13
timestamp 1635444444
transform 1 0 2300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_21
timestamp 1635444444
transform 1 0 3036 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _312_
timestamp 1635444444
transform -1 0 3036 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1635444444
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1635444444
transform 1 0 4048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1635444444
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _288_
timestamp 1635444444
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1635444444
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1635444444
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1635444444
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1635444444
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1635444444
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1635444444
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _292_
timestamp 1635444444
transform -1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_91
timestamp 1635444444
transform 1 0 9476 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_99
timestamp 1635444444
transform 1 0 10212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1635444444
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1635444444
transform -1 0 10856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1635444444
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1635444444
transform 1 0 1380 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1635444444
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_21
timestamp 1635444444
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _311_
timestamp 1635444444
transform -1 0 3036 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_33
timestamp 1635444444
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1635444444
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1635444444
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1635444444
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1635444444
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1635444444
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1635444444
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_93
timestamp 1635444444
transform 1 0 9660 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_99
timestamp 1635444444
transform 1 0 10212 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _291_
timestamp 1635444444
transform 1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1635444444
transform -1 0 10856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1635444444
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1635444444
transform 1 0 1380 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_18_13
timestamp 1635444444
transform 1 0 2300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1635444444
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _313_
timestamp 1635444444
transform -1 0 3036 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1635444444
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1635444444
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1635444444
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1635444444
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1635444444
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1635444444
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1635444444
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1635444444
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1635444444
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1635444444
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1635444444
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1635444444
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1635444444
transform 1 0 9844 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1635444444
transform -1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1635444444
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1635444444
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1635444444
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1635444444
transform 1 0 1380 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1635444444
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1635444444
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_17
timestamp 1635444444
transform 1 0 2668 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1635444444
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1635444444
transform 1 0 2668 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1635444444
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1635444444
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1635444444
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_37
timestamp 1635444444
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1635444444
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _216_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 4508 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1635444444
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1635444444
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_49
timestamp 1635444444
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1635444444
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1635444444
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_61
timestamp 1635444444
transform 1 0 6716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1635444444
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1635444444
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1635444444
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_81
timestamp 1635444444
transform 1 0 8556 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp 1635444444
transform 1 0 9108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1635444444
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1635444444
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1635444444
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _296_
timestamp 1635444444
transform -1 0 9476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1635444444
transform 1 0 9476 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_99
timestamp 1635444444
transform 1 0 10212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1635444444
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99
timestamp 1635444444
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1635444444
transform 1 0 9844 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1635444444
transform 1 0 9844 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1635444444
transform -1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1635444444
transform -1 0 10856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_11
timestamp 1635444444
transform 1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1635444444
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1635444444
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1635444444
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1635444444
transform 1 0 2760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_25
timestamp 1635444444
transform 1 0 3404 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1635444444
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _289_
timestamp 1635444444
transform -1 0 3404 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_32
timestamp 1635444444
transform 1 0 4048 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _290_
timestamp 1635444444
transform -1 0 4048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1635444444
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1635444444
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1635444444
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1635444444
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1635444444
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1635444444
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1635444444
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1635444444
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1635444444
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_93
timestamp 1635444444
transform 1 0 9660 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1635444444
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_3
timestamp 1635444444
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1635444444
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2392 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_22_14
timestamp 1635444444
transform 1 0 2392 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_20
timestamp 1635444444
transform 1 0 2944 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1635444444
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _228_
timestamp 1635444444
transform -1 0 3312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1635444444
transform 1 0 4048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1635444444
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1635444444
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1635444444
transform 1 0 4416 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_39
timestamp 1635444444
transform 1 0 4692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_51
timestamp 1635444444
transform 1 0 5796 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1635444444
transform 1 0 6900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_75
timestamp 1635444444
transform 1 0 8004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1635444444
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1635444444
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1635444444
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1635444444
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_99
timestamp 1635444444
transform 1 0 10212 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1635444444
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1635444444
transform -1 0 10856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_9
timestamp 1635444444
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1635444444
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 1932 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_18
timestamp 1635444444
transform 1 0 2760 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _271_
timestamp 1635444444
transform -1 0 2760 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _272_
timestamp 1635444444
transform 1 0 3128 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1635444444
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1635444444
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1635444444
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1635444444
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1635444444
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1635444444
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1635444444
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_81
timestamp 1635444444
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1635444444
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1635444444
transform -1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1635444444
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1635444444
transform 1 0 10212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1635444444
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1635444444
transform -1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_6
timestamp 1635444444
transform 1 0 1656 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1635444444
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _083_
timestamp 1635444444
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1635444444
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _089_
timestamp 1635444444
transform 1 0 2392 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1635444444
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1635444444
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1635444444
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1635444444
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1635444444
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1635444444
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1635444444
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1635444444
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1635444444
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1635444444
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1635444444
transform 1 0 9660 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1635444444
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _298_
timestamp 1635444444
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1635444444
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_10
timestamp 1635444444
transform 1 0 2024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1635444444
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1635444444
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _085_
timestamp 1635444444
transform 1 0 1472 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_17
timestamp 1635444444
transform 1 0 2668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_24
timestamp 1635444444
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1635444444
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1635444444
transform 1 0 3036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_36
timestamp 1635444444
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1635444444
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1635444444
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1635444444
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1635444444
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_81
timestamp 1635444444
transform 1 0 8556 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_87
timestamp 1635444444
transform 1 0 9108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _299_
timestamp 1635444444
transform -1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_91
timestamp 1635444444
transform 1 0 9476 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_99
timestamp 1635444444
transform 1 0 10212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1635444444
transform 1 0 9844 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1635444444
transform -1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_6
timestamp 1635444444
transform 1 0 1656 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1635444444
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1635444444
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1635444444
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1635444444
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1635444444
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1635444444
transform 1 0 2024 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_14
timestamp 1635444444
transform 1 0 2392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_22
timestamp 1635444444
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_13
timestamp 1635444444
transform 1 0 2300 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_20
timestamp 1635444444
transform 1 0 2944 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_1  _090_
timestamp 1635444444
transform -1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1635444444
transform 1 0 2668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1635444444
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1635444444
transform 1 0 4048 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1635444444
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1635444444
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1635444444
transform 1 0 5152 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1635444444
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1635444444
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1635444444
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1635444444
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1635444444
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1635444444
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1635444444
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1635444444
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1635444444
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1635444444
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _297_
timestamp 1635444444
transform -1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_91
timestamp 1635444444
transform 1 0 9476 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1635444444
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1635444444
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_99
timestamp 1635444444
transform 1 0 10212 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1635444444
transform 1 0 9844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1635444444
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1635444444
transform -1 0 10856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1635444444
transform -1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1635444444
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_9
timestamp 1635444444
transform 1 0 1932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1635444444
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1635444444
transform 1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_20
timestamp 1635444444
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _088_
timestamp 1635444444
transform 1 0 2484 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1635444444
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1635444444
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1635444444
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1635444444
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1635444444
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1635444444
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1635444444
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_85
timestamp 1635444444
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1635444444
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_102
timestamp 1635444444
transform 1 0 10488 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1635444444
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1635444444
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _300_
timestamp 1635444444
transform 1 0 9844 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1635444444
transform -1 0 10856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_6
timestamp 1635444444
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1635444444
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1635444444
transform -1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1635444444
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1635444444
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_20
timestamp 1635444444
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1635444444
transform 1 0 2668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1635444444
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1635444444
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1635444444
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1635444444
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1635444444
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1635444444
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1635444444
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_99
timestamp 1635444444
transform 1 0 10212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1635444444
transform 1 0 9844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1635444444
transform -1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_10
timestamp 1635444444
transform 1 0 2024 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1635444444
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1635444444
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1635444444
transform -1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_17
timestamp 1635444444
transform 1 0 2668 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1635444444
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1635444444
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1635444444
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1635444444
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1635444444
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1635444444
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1635444444
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1635444444
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1635444444
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1635444444
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1635444444
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1635444444
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _301_
timestamp 1635444444
transform -1 0 9476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1635444444
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_99
timestamp 1635444444
transform 1 0 10212 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1635444444
transform 1 0 9844 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1635444444
transform -1 0 10856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_6
timestamp 1635444444
transform 1 0 1656 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1635444444
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1635444444
transform -1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1635444444
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_15
timestamp 1635444444
transform 1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_22
timestamp 1635444444
transform 1 0 3128 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1635444444
transform 1 0 2852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_34
timestamp 1635444444
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_46
timestamp 1635444444
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1635444444
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1635444444
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1635444444
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1635444444
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1635444444
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_93
timestamp 1635444444
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1635444444
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _302_
timestamp 1635444444
transform 1 0 9936 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1635444444
transform -1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_11
timestamp 1635444444
transform 1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1635444444
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1635444444
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1635444444
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1635444444
transform -1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 1635444444
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1635444444
transform -1 0 2760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1635444444
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1635444444
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_37
timestamp 1635444444
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1635444444
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _227_
timestamp 1635444444
transform -1 0 4508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_49
timestamp 1635444444
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_61
timestamp 1635444444
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1635444444
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1635444444
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1635444444
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1635444444
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1635444444
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1635444444
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1635444444
transform 1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1635444444
transform -1 0 10856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1635444444
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_7
timestamp 1635444444
transform 1 0 1748 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_11
timestamp 1635444444
transform 1 0 2116 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1635444444
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_7
timestamp 1635444444
transform 1 0 1748 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1635444444
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1635444444
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1635444444
transform -1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1635444444
transform -1 0 2116 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_19
timestamp 1635444444
transform 1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1635444444
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2484 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1635444444
transform -1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input128
timestamp 1635444444
transform 1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_26
timestamp 1635444444
transform 1 0 3496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_33
timestamp 1635444444
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1635444444
transform 1 0 4048 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1635444444
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1635444444
transform 1 0 3864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input130
timestamp 1635444444
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1635444444
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1635444444
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1635444444
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1635444444
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1635444444
transform 1 0 6256 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1635444444
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_69
timestamp 1635444444
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1635444444
transform 1 0 7360 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_81
timestamp 1635444444
transform 1 0 8556 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_87
timestamp 1635444444
transform 1 0 9108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1635444444
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1635444444
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1635444444
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _303_
timestamp 1635444444
transform -1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1635444444
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_99
timestamp 1635444444
transform 1 0 10212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1635444444
transform 1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1635444444
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1635444444
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1635444444
transform 1 0 9844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1635444444
transform -1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1635444444
transform -1 0 10856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_10
timestamp 1635444444
transform 1 0 2024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1635444444
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1635444444
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1635444444
transform -1 0 2024 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_14
timestamp 1635444444
transform 1 0 2392 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_24
timestamp 1635444444
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_4  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 2484 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_35_31
timestamp 1635444444
transform 1 0 3956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1635444444
transform 1 0 3680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_43
timestamp 1635444444
transform 1 0 5060 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1635444444
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1635444444
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1635444444
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_69
timestamp 1635444444
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_81
timestamp 1635444444
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_101
timestamp 1635444444
transform 1 0 10396 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_93
timestamp 1635444444
transform 1 0 9660 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1635444444
transform -1 0 10856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1635444444
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1635444444
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _114_
timestamp 1635444444
transform -1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_13
timestamp 1635444444
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_20
timestamp 1635444444
transform 1 0 2944 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1635444444
transform 1 0 2668 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1635444444
transform 1 0 4048 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1635444444
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1635444444
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1635444444
transform 1 0 5152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1635444444
transform 1 0 6256 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1635444444
transform 1 0 7360 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1635444444
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1635444444
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1635444444
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1635444444
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_99
timestamp 1635444444
transform 1 0 10212 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1635444444
transform 1 0 9844 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1635444444
transform -1 0 10856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1635444444
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_9
timestamp 1635444444
transform 1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1635444444
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _118_
timestamp 1635444444
transform -1 0 1932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_16
timestamp 1635444444
transform 1 0 2576 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_23
timestamp 1635444444
transform 1 0 3220 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1635444444
transform -1 0 2576 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1635444444
transform 1 0 2944 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_35
timestamp 1635444444
transform 1 0 4324 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_47
timestamp 1635444444
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1635444444
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1635444444
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1635444444
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1635444444
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1635444444
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1635444444
transform 1 0 9660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_99
timestamp 1635444444
transform 1 0 10212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1635444444
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1635444444
transform -1 0 10856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1635444444
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1635444444
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _120_
timestamp 1635444444
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _124_
timestamp 1635444444
transform 1 0 2116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1635444444
transform 1 0 2484 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1635444444
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _126_
timestamp 1635444444
transform 1 0 2852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1635444444
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1635444444
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1635444444
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1635444444
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1635444444
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1635444444
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1635444444
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1635444444
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1635444444
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1635444444
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _304_
timestamp 1635444444
transform -1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_92
timestamp 1635444444
transform 1 0 9568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_99
timestamp 1635444444
transform 1 0 10212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 9936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1635444444
transform -1 0 10856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_6
timestamp 1635444444
transform 1 0 1656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_6
timestamp 1635444444
transform 1 0 1656 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1635444444
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1635444444
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _129_
timestamp 1635444444
transform -1 0 2576 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _131_
timestamp 1635444444
transform 1 0 2208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1635444444
transform -1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1635444444
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_16
timestamp 1635444444
transform 1 0 2576 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_16
timestamp 1635444444
transform 1 0 2576 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_23
timestamp 1635444444
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1635444444
transform 1 0 2944 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_28
timestamp 1635444444
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1635444444
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1635444444
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1635444444
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_40
timestamp 1635444444
transform 1 0 4784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1635444444
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1635444444
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1635444444
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1635444444
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1635444444
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1635444444
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1635444444
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1635444444
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1635444444
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1635444444
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1635444444
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1635444444
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_93
timestamp 1635444444
transform 1 0 9660 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1635444444
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1635444444
transform 1 0 9660 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_99
timestamp 1635444444
transform 1 0 10212 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _276_
timestamp 1635444444
transform 1 0 9936 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1635444444
transform 1 0 9844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1635444444
transform -1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1635444444
transform -1 0 10856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_6
timestamp 1635444444
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1635444444
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _133_
timestamp 1635444444
transform -1 0 2392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1635444444
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_14
timestamp 1635444444
transform 1 0 2392 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _215_
timestamp 1635444444
transform 1 0 2944 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_26
timestamp 1635444444
transform 1 0 3496 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_38
timestamp 1635444444
transform 1 0 4600 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_50
timestamp 1635444444
transform 1 0 5704 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1635444444
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1635444444
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1635444444
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1635444444
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_93
timestamp 1635444444
transform 1 0 9660 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1635444444
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _277_
timestamp 1635444444
transform 1 0 9936 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1635444444
transform -1 0 10856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1635444444
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_9
timestamp 1635444444
transform 1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1635444444
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _135_
timestamp 1635444444
transform -1 0 1932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_17
timestamp 1635444444
transform 1 0 2668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1635444444
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _137_
timestamp 1635444444
transform 1 0 2300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1635444444
transform 1 0 3036 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1635444444
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1635444444
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1635444444
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1635444444
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1635444444
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1635444444
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1635444444
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1635444444
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1635444444
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_93
timestamp 1635444444
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_99
timestamp 1635444444
transform 1 0 10212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _278_
timestamp 1635444444
transform 1 0 9936 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1635444444
transform -1 0 10856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_12
timestamp 1635444444
transform 1 0 2208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_3
timestamp 1635444444
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_7
timestamp 1635444444
transform 1 0 1748 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1635444444
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _140_
timestamp 1635444444
transform 1 0 1840 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_19
timestamp 1635444444
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1635444444
transform 1 0 2576 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_31
timestamp 1635444444
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_43
timestamp 1635444444
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1635444444
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1635444444
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1635444444
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1635444444
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1635444444
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_101
timestamp 1635444444
transform 1 0 10396 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_93
timestamp 1635444444
transform 1 0 9660 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1635444444
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_6
timestamp 1635444444
transform 1 0 1656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1635444444
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1635444444
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1635444444
transform -1 0 2300 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_13
timestamp 1635444444
transform 1 0 2300 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_19
timestamp 1635444444
transform 1 0 2852 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1635444444
transform 1 0 3220 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _232_
timestamp 1635444444
transform -1 0 3220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1635444444
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1635444444
transform 1 0 4048 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1635444444
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1635444444
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1635444444
transform 1 0 5152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_56
timestamp 1635444444
transform 1 0 6256 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1635444444
transform 1 0 7360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1635444444
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1635444444
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1635444444
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_97
timestamp 1635444444
transform 1 0 10028 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1635444444
transform -1 0 10856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1635444444
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_9
timestamp 1635444444
transform 1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1635444444
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _142_
timestamp 1635444444
transform -1 0 1932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_18
timestamp 1635444444
transform 1 0 2760 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _093_
timestamp 1635444444
transform -1 0 3496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _096_
timestamp 1635444444
transform -1 0 2760 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_45_26
timestamp 1635444444
transform 1 0 3496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_33
timestamp 1635444444
transform 1 0 4140 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _231_
timestamp 1635444444
transform -1 0 4140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1635444444
transform 1 0 4508 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_40
timestamp 1635444444
transform 1 0 4784 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1635444444
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1635444444
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1635444444
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1635444444
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1635444444
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_93
timestamp 1635444444
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1635444444
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _273_
timestamp 1635444444
transform -1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1635444444
transform -1 0 10856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1635444444
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_3
timestamp 1635444444
transform 1 0 1380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_8
timestamp 1635444444
transform 1 0 1840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1635444444
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1635444444
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _094_
timestamp 1635444444
transform -1 0 2668 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _100_
timestamp 1635444444
transform 1 0 2024 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_2  _148_
timestamp 1635444444
transform -1 0 1840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1635444444
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1635444444
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1635444444
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_17
timestamp 1635444444
transform 1 0 2668 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_25
timestamp 1635444444
transform 1 0 3404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1635444444
transform -1 0 3404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _230_
timestamp 1635444444
transform -1 0 3312 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1635444444
transform 1 0 4048 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_32
timestamp 1635444444
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1635444444
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp 1635444444
transform -1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input116
timestamp 1635444444
transform 1 0 3772 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1635444444
transform 1 0 5152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_44
timestamp 1635444444
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1635444444
transform 1 0 6256 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1635444444
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1635444444
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1635444444
transform 1 0 7360 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1635444444
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1635444444
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1635444444
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1635444444
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1635444444
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1635444444
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_99
timestamp 1635444444
transform 1 0 10212 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_101
timestamp 1635444444
transform 1 0 10396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_93
timestamp 1635444444
transform 1 0 9660 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _274_
timestamp 1635444444
transform -1 0 10212 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1635444444
transform -1 0 10856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1635444444
transform -1 0 10856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_11
timestamp 1635444444
transform 1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_3
timestamp 1635444444
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1635444444
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _144_
timestamp 1635444444
transform -1 0 2116 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 1635444444
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _146_
timestamp 1635444444
transform -1 0 2852 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1635444444
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1635444444
transform 1 0 4048 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1635444444
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1635444444
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1635444444
transform 1 0 5152 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1635444444
transform 1 0 6256 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1635444444
transform 1 0 7360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1635444444
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1635444444
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1635444444
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_97
timestamp 1635444444
transform 1 0 10028 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1635444444
transform -1 0 10856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_3
timestamp 1635444444
transform 1 0 1380 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1635444444
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _098_
timestamp 1635444444
transform 1 0 1932 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_49_14
timestamp 1635444444
transform 1 0 2392 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_23
timestamp 1635444444
transform 1 0 3220 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _102_
timestamp 1635444444
transform -1 0 3220 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_49_30
timestamp 1635444444
transform 1 0 3864 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1635444444
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_42
timestamp 1635444444
transform 1 0 4968 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1635444444
transform 1 0 6072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1635444444
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1635444444
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1635444444
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1635444444
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_93
timestamp 1635444444
transform 1 0 9660 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_99
timestamp 1635444444
transform 1 0 10212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _279_
timestamp 1635444444
transform 1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1635444444
transform -1 0 10856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_3
timestamp 1635444444
transform 1 0 1380 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_8
timestamp 1635444444
transform 1 0 1840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1635444444
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _162_
timestamp 1635444444
transform -1 0 1840 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1635444444
transform 1 0 2208 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1635444444
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_22
timestamp 1635444444
transform 1 0 3128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1635444444
transform 1 0 2852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1635444444
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1635444444
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1635444444
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1635444444
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1635444444
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1635444444
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1635444444
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1635444444
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1635444444
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_97
timestamp 1635444444
transform 1 0 10028 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1635444444
transform -1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_3
timestamp 1635444444
transform 1 0 1380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_7
timestamp 1635444444
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1635444444
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1635444444
transform -1 0 1748 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input121
timestamp 1635444444
transform -1 0 2392 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_14
timestamp 1635444444
transform 1 0 2392 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_21
timestamp 1635444444
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1635444444
transform 1 0 2760 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_33
timestamp 1635444444
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_45
timestamp 1635444444
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1635444444
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1635444444
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1635444444
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1635444444
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1635444444
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_93
timestamp 1635444444
transform 1 0 9660 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_99
timestamp 1635444444
transform 1 0 10212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1635444444
transform 1 0 9844 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1635444444
transform -1 0 10856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_7
timestamp 1635444444
transform 1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_3
timestamp 1635444444
transform 1 0 1380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_8
timestamp 1635444444
transform 1 0 1840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1635444444
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1635444444
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _153_
timestamp 1635444444
transform -1 0 1840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1635444444
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1635444444
transform -1 0 1748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output262
timestamp 1635444444
transform 1 0 2208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_14
timestamp 1635444444
transform 1 0 2392 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_16
timestamp 1635444444
transform 1 0 2576 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_26
timestamp 1635444444
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1635444444
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_28
timestamp 1635444444
transform 1 0 3680 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1635444444
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1635444444
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_40
timestamp 1635444444
transform 1 0 4784 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1635444444
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1635444444
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1635444444
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1635444444
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1635444444
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1635444444
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1635444444
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1635444444
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_85
timestamp 1635444444
transform 1 0 8924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1635444444
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1635444444
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_93
timestamp 1635444444
transform 1 0 9660 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_99
timestamp 1635444444
transform 1 0 10212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1635444444
transform 1 0 9660 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_99
timestamp 1635444444
transform 1 0 10212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _280_
timestamp 1635444444
transform 1 0 9936 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1635444444
transform 1 0 9844 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1635444444
transform -1 0 10856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1635444444
transform -1 0 10856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1635444444
transform 1 0 1380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_8
timestamp 1635444444
transform 1 0 1840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1635444444
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _155_
timestamp 1635444444
transform -1 0 1840 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1635444444
transform 1 0 2208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_16
timestamp 1635444444
transform 1 0 2576 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1635444444
transform 1 0 4048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1635444444
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1635444444
transform -1 0 4048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1635444444
transform 1 0 5152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1635444444
transform 1 0 6256 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1635444444
transform 1 0 7360 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1635444444
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1635444444
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1635444444
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1635444444
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1635444444
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1635444444
transform 1 0 9844 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1635444444
transform -1 0 10856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_6
timestamp 1635444444
transform 1 0 1656 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1635444444
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _105_
timestamp 1635444444
transform 1 0 2024 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _268_
timestamp 1635444444
transform -1 0 1656 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_15
timestamp 1635444444
transform 1 0 2484 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _236_
timestamp 1635444444
transform -1 0 3496 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_26
timestamp 1635444444
transform 1 0 3496 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_38
timestamp 1635444444
transform 1 0 4600 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_50
timestamp 1635444444
transform 1 0 5704 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1635444444
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1635444444
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1635444444
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1635444444
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_93
timestamp 1635444444
transform 1 0 9660 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_99
timestamp 1635444444
transform 1 0 10212 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1635444444
transform 1 0 9844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1635444444
transform -1 0 10856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_7
timestamp 1635444444
transform 1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1635444444
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output276
timestamp 1635444444
transform -1 0 1748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1635444444
transform 1 0 2116 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_15
timestamp 1635444444
transform 1 0 2484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_22
timestamp 1635444444
transform 1 0 3128 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _267_
timestamp 1635444444
transform 1 0 2852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1635444444
transform 1 0 4048 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1635444444
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1635444444
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1635444444
transform 1 0 5152 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1635444444
transform 1 0 6256 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1635444444
transform 1 0 7360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1635444444
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1635444444
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1635444444
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_97
timestamp 1635444444
transform 1 0 10028 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1635444444
transform -1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_11
timestamp 1635444444
transform 1 0 2116 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_7
timestamp 1635444444
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1635444444
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _107_
timestamp 1635444444
transform -1 0 2668 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output277
timestamp 1635444444
transform -1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_17
timestamp 1635444444
transform 1 0 2668 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_24
timestamp 1635444444
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _237_
timestamp 1635444444
transform -1 0 3312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_36
timestamp 1635444444
transform 1 0 4416 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_48
timestamp 1635444444
transform 1 0 5520 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1635444444
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1635444444
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1635444444
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1635444444
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_93
timestamp 1635444444
transform 1 0 9660 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_99
timestamp 1635444444
transform 1 0 10212 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1635444444
transform 1 0 9844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1635444444
transform -1 0 10856 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_7
timestamp 1635444444
transform 1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1635444444
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1635444444
transform -1 0 1748 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output280
timestamp 1635444444
transform 1 0 2116 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_15
timestamp 1635444444
transform 1 0 2484 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_23
timestamp 1635444444
transform 1 0 3220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1635444444
transform 1 0 2852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1635444444
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1635444444
transform 1 0 4048 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1635444444
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _239_
timestamp 1635444444
transform -1 0 4048 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1635444444
transform 1 0 5152 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1635444444
transform 1 0 6256 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1635444444
transform 1 0 7360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1635444444
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_85
timestamp 1635444444
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1635444444
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1635444444
transform 1 0 9660 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_99
timestamp 1635444444
transform 1 0 10212 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1635444444
transform 1 0 9844 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1635444444
transform -1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1635444444
transform -1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _159_
timestamp 1635444444
transform -1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1635444444
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1635444444
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1635444444
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_11
timestamp 1635444444
transform 1 0 2116 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_7
timestamp 1635444444
transform 1 0 1748 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_11
timestamp 1635444444
transform 1 0 2116 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _111_
timestamp 1635444444
transform 1 0 2208 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _109_
timestamp 1635444444
transform 1 0 2208 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_59_17
timestamp 1635444444
transform 1 0 2668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_25
timestamp 1635444444
transform 1 0 3404 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_17
timestamp 1635444444
transform 1 0 2668 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_24
timestamp 1635444444
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _238_
timestamp 1635444444
transform -1 0 3312 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1635444444
transform 1 0 3036 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_37
timestamp 1635444444
transform 1 0 4508 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1635444444
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1635444444
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1635444444
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1635444444
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1635444444
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1635444444
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1635444444
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1635444444
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1635444444
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1635444444
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1635444444
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1635444444
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1635444444
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1635444444
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1635444444
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_101
timestamp 1635444444
transform 1 0 10396 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_93
timestamp 1635444444
transform 1 0 9660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_93
timestamp 1635444444
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_99
timestamp 1635444444
transform 1 0 10212 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1635444444
transform 1 0 9844 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1635444444
transform -1 0 10856 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1635444444
transform -1 0 10856 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_3
timestamp 1635444444
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_9
timestamp 1635444444
transform 1 0 1932 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1635444444
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _163_
timestamp 1635444444
transform -1 0 1932 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_61_13
timestamp 1635444444
transform 1 0 2300 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_19
timestamp 1635444444
transform 1 0 2852 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _113_
timestamp 1635444444
transform -1 0 2852 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _234_
timestamp 1635444444
transform 1 0 3404 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_61_35
timestamp 1635444444
transform 1 0 4324 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_47
timestamp 1635444444
transform 1 0 5428 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1635444444
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1635444444
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1635444444
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1635444444
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1635444444
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_93
timestamp 1635444444
transform 1 0 9660 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_99
timestamp 1635444444
transform 1 0 10212 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1635444444
transform 1 0 9844 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1635444444
transform -1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1635444444
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1635444444
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1635444444
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1635444444
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1635444444
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1635444444
transform 1 0 4048 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1635444444
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _241_
timestamp 1635444444
transform -1 0 4048 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1635444444
transform 1 0 5152 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1635444444
transform 1 0 6256 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1635444444
transform 1 0 7360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1635444444
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_85
timestamp 1635444444
transform 1 0 8924 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1635444444
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1635444444
transform 1 0 9660 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_99
timestamp 1635444444
transform 1 0 10212 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1635444444
transform 1 0 9844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1635444444
transform -1 0 10856 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_7
timestamp 1635444444
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1635444444
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1635444444
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1635444444
transform -1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1635444444
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_23
timestamp 1635444444
transform 1 0 3220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1635444444
transform 1 0 2852 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_30
timestamp 1635444444
transform 1 0 3864 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _242_
timestamp 1635444444
transform -1 0 3864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_42
timestamp 1635444444
transform 1 0 4968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1635444444
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1635444444
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1635444444
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1635444444
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1635444444
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_101
timestamp 1635444444
transform 1 0 10396 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_93
timestamp 1635444444
transform 1 0 9660 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1635444444
transform -1 0 10856 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_8
timestamp 1635444444
transform 1 0 1840 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1635444444
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _161_
timestamp 1635444444
transform 1 0 1380 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1635444444
transform -1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_16
timestamp 1635444444
transform 1 0 2576 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_23
timestamp 1635444444
transform 1 0 3220 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1635444444
transform 1 0 2944 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1635444444
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1635444444
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1635444444
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1635444444
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1635444444
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1635444444
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1635444444
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1635444444
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1635444444
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1635444444
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1635444444
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_99
timestamp 1635444444
transform 1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1635444444
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1635444444
transform -1 0 10856 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_11
timestamp 1635444444
transform 1 0 2116 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_7
timestamp 1635444444
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1635444444
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _149_
timestamp 1635444444
transform -1 0 2576 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1635444444
transform -1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_16
timestamp 1635444444
transform 1 0 2576 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_28
timestamp 1635444444
transform 1 0 3680 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_40
timestamp 1635444444
transform 1 0 4784 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_52
timestamp 1635444444
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1635444444
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1635444444
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1635444444
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1635444444
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_93
timestamp 1635444444
transform 1 0 9660 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_99
timestamp 1635444444
transform 1 0 10212 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1635444444
transform 1 0 9844 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1635444444
transform -1 0 10856 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_3
timestamp 1635444444
transform 1 0 1380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_9
timestamp 1635444444
transform 1 0 1932 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_11
timestamp 1635444444
transform 1 0 2116 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_3
timestamp 1635444444
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1635444444
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1635444444
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _121_
timestamp 1635444444
transform -1 0 2116 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1635444444
transform -1 0 2392 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_14
timestamp 1635444444
transform 1 0 2392 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_22
timestamp 1635444444
transform 1 0 3128 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_23
timestamp 1635444444
transform 1 0 3220 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1635444444
transform -1 0 3128 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _233_
timestamp 1635444444
transform 1 0 2852 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1635444444
transform 1 0 4048 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_30
timestamp 1635444444
transform 1 0 3864 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_37
timestamp 1635444444
transform 1 0 4508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1635444444
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _243_
timestamp 1635444444
transform -1 0 3864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1635444444
transform -1 0 4508 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _248_
timestamp 1635444444
transform -1 0 4048 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1635444444
transform 1 0 5152 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_49
timestamp 1635444444
transform 1 0 5612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1635444444
transform 1 0 6256 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1635444444
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1635444444
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1635444444
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1635444444
transform 1 0 7360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1635444444
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1635444444
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1635444444
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1635444444
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1635444444
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_97
timestamp 1635444444
transform 1 0 10028 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_93
timestamp 1635444444
transform 1 0 9660 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_99
timestamp 1635444444
transform 1 0 10212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1635444444
transform 1 0 9844 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1635444444
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1635444444
transform -1 0 10856 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_7
timestamp 1635444444
transform 1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1635444444
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output259
timestamp 1635444444
transform -1 0 1748 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output260
timestamp 1635444444
transform -1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_15
timestamp 1635444444
transform 1 0 2484 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_23
timestamp 1635444444
transform 1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output261
timestamp 1635444444
transform -1 0 3220 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1635444444
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_32
timestamp 1635444444
transform 1 0 4048 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1635444444
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _117_
timestamp 1635444444
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 1635444444
transform -1 0 4692 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_39
timestamp 1635444444
transform 1 0 4692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_51
timestamp 1635444444
transform 1 0 5796 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_63
timestamp 1635444444
transform 1 0 6900 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_75
timestamp 1635444444
transform 1 0 8004 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1635444444
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_85
timestamp 1635444444
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1635444444
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_93
timestamp 1635444444
transform 1 0 9660 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_99
timestamp 1635444444
transform 1 0 10212 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1635444444
transform 1 0 9844 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1635444444
transform -1 0 10856 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_3
timestamp 1635444444
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_7
timestamp 1635444444
transform 1 0 1748 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1635444444
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _125_
timestamp 1635444444
transform -1 0 2300 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_69_13
timestamp 1635444444
transform 1 0 2300 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_21
timestamp 1635444444
transform 1 0 3036 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1635444444
transform 1 0 2668 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _123_
timestamp 1635444444
transform 1 0 3404 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_28
timestamp 1635444444
transform 1 0 3680 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_35
timestamp 1635444444
transform 1 0 4324 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _245_
timestamp 1635444444
transform -1 0 4324 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_47
timestamp 1635444444
transform 1 0 5428 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1635444444
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1635444444
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1635444444
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1635444444
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1635444444
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_93
timestamp 1635444444
transform 1 0 9660 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_99
timestamp 1635444444
transform 1 0 10212 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1635444444
transform 1 0 9844 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1635444444
transform -1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_7
timestamp 1635444444
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1635444444
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output263
timestamp 1635444444
transform -1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1635444444
transform 1 0 2116 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_15
timestamp 1635444444
transform 1 0 2484 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_23
timestamp 1635444444
transform 1 0 3220 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1635444444
transform 1 0 2852 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1635444444
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_32
timestamp 1635444444
transform 1 0 4048 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1635444444
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _119_
timestamp 1635444444
transform 1 0 3772 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_44
timestamp 1635444444
transform 1 0 5152 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_56
timestamp 1635444444
transform 1 0 6256 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_68
timestamp 1635444444
transform 1 0 7360 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_80
timestamp 1635444444
transform 1 0 8464 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1635444444
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1635444444
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_97
timestamp 1635444444
transform 1 0 10028 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1635444444
transform -1 0 10856 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_3
timestamp 1635444444
transform 1 0 1380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_9
timestamp 1635444444
transform 1 0 1932 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1635444444
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _150_
timestamp 1635444444
transform 1 0 1472 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_71_17
timestamp 1635444444
transform 1 0 2668 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1635444444
transform -1 0 2668 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_29
timestamp 1635444444
transform 1 0 3772 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_41
timestamp 1635444444
transform 1 0 4876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1635444444
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1635444444
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1635444444
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1635444444
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1635444444
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_93
timestamp 1635444444
transform 1 0 9660 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_99
timestamp 1635444444
transform 1 0 10212 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1635444444
transform 1 0 9844 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1635444444
transform -1 0 10856 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_7
timestamp 1635444444
transform 1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_7
timestamp 1635444444
transform 1 0 1748 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1635444444
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1635444444
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _315_
timestamp 1635444444
transform 1 0 2116 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1635444444
transform -1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output268
timestamp 1635444444
transform -1 0 1748 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_14
timestamp 1635444444
transform 1 0 2392 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_19
timestamp 1635444444
transform 1 0 2852 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_23
timestamp 1635444444
transform 1 0 3220 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _240_
timestamp 1635444444
transform 1 0 3312 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 1635444444
transform 1 0 3496 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_29
timestamp 1635444444
transform 1 0 3772 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_33
timestamp 1635444444
transform 1 0 4140 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_28
timestamp 1635444444
transform 1 0 3680 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_36
timestamp 1635444444
transform 1 0 4416 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1635444444
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _246_
timestamp 1635444444
transform 1 0 4048 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1635444444
transform -1 0 4140 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_45
timestamp 1635444444
transform 1 0 5244 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_48
timestamp 1635444444
transform 1 0 5520 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_57
timestamp 1635444444
transform 1 0 6348 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1635444444
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1635444444
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_69
timestamp 1635444444
transform 1 0 7452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1635444444
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_81
timestamp 1635444444
transform 1 0 8556 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1635444444
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1635444444
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1635444444
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_93
timestamp 1635444444
transform 1 0 9660 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_99
timestamp 1635444444
transform 1 0 10212 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_101
timestamp 1635444444
transform 1 0 10396 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_93
timestamp 1635444444
transform 1 0 9660 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1635444444
transform 1 0 9844 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1635444444
transform -1 0 10856 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1635444444
transform -1 0 10856 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_7
timestamp 1635444444
transform 1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1635444444
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1635444444
transform -1 0 1748 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output271
timestamp 1635444444
transform -1 0 2484 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1635444444
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1635444444
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1635444444
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1635444444
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1635444444
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1635444444
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1635444444
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1635444444
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1635444444
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_85
timestamp 1635444444
transform 1 0 8924 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1635444444
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_93
timestamp 1635444444
transform 1 0 9660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_99
timestamp 1635444444
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1635444444
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1635444444
transform -1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_7
timestamp 1635444444
transform 1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1635444444
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _132_
timestamp 1635444444
transform 1 0 2116 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output270
timestamp 1635444444
transform -1 0 1748 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_14
timestamp 1635444444
transform 1 0 2392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1635444444
transform 1 0 2760 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_75_28
timestamp 1635444444
transform 1 0 3680 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_40
timestamp 1635444444
transform 1 0 4784 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_52
timestamp 1635444444
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1635444444
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1635444444
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1635444444
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1635444444
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_93
timestamp 1635444444
transform 1 0 9660 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_99
timestamp 1635444444
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1635444444
transform 1 0 9844 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1635444444
transform -1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_7
timestamp 1635444444
transform 1 0 1748 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1635444444
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1635444444
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output272
timestamp 1635444444
transform -1 0 2484 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_15
timestamp 1635444444
transform 1 0 2484 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_23
timestamp 1635444444
transform 1 0 3220 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output274
timestamp 1635444444
transform 1 0 2852 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1635444444
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_29
timestamp 1635444444
transform 1 0 3772 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_37
timestamp 1635444444
transform 1 0 4508 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1635444444
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _258_
timestamp 1635444444
transform 1 0 4140 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1635444444
transform 1 0 5152 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _250_
timestamp 1635444444
transform -1 0 5152 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_56
timestamp 1635444444
transform 1 0 6256 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_68
timestamp 1635444444
transform 1 0 7360 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_80
timestamp 1635444444
transform 1 0 8464 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_85
timestamp 1635444444
transform 1 0 8924 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1635444444
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_93
timestamp 1635444444
transform 1 0 9660 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_99
timestamp 1635444444
transform 1 0 10212 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1635444444
transform 1 0 9844 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1635444444
transform -1 0 10856 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_77_3
timestamp 1635444444
transform 1 0 1380 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_9
timestamp 1635444444
transform 1 0 1932 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1635444444
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _152_
timestamp 1635444444
transform 1 0 1472 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_77_17
timestamp 1635444444
transform 1 0 2668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_24
timestamp 1635444444
transform 1 0 3312 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _130_
timestamp 1635444444
transform 1 0 3036 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output275
timestamp 1635444444
transform 1 0 2300 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_31
timestamp 1635444444
transform 1 0 3956 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_38
timestamp 1635444444
transform 1 0 4600 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _134_
timestamp 1635444444
transform 1 0 3680 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _261_
timestamp 1635444444
transform -1 0 4600 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_50
timestamp 1635444444
transform 1 0 5704 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1635444444
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1635444444
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1635444444
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1635444444
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_101
timestamp 1635444444
transform 1 0 10396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1635444444
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1635444444
transform -1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_3
timestamp 1635444444
transform 1 0 1380 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_9
timestamp 1635444444
transform 1 0 1932 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1635444444
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _156_
timestamp 1635444444
transform -1 0 1932 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_78_17
timestamp 1635444444
transform 1 0 2668 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_24
timestamp 1635444444
transform 1 0 3312 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _253_
timestamp 1635444444
transform -1 0 3312 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1635444444
transform -1 0 2668 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1635444444
transform 1 0 4048 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1635444444
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _251_
timestamp 1635444444
transform -1 0 4048 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_44
timestamp 1635444444
transform 1 0 5152 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_56
timestamp 1635444444
transform 1 0 6256 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_68
timestamp 1635444444
transform 1 0 7360 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1635444444
transform 1 0 8464 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_78_85
timestamp 1635444444
transform 1 0 8924 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1635444444
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_93
timestamp 1635444444
transform 1 0 9660 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_99
timestamp 1635444444
transform 1 0 10212 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1635444444
transform 1 0 9844 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1635444444
transform -1 0 10856 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_7
timestamp 1635444444
transform 1 0 1748 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_11
timestamp 1635444444
transform 1 0 2116 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_80_3
timestamp 1635444444
transform 1 0 1380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1635444444
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1635444444
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _158_
timestamp 1635444444
transform -1 0 2116 0 1 45696
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1635444444
transform -1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_19
timestamp 1635444444
transform 1 0 2852 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_80_19
timestamp 1635444444
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _252_
timestamp 1635444444
transform 1 0 3404 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1635444444
transform 1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_35
timestamp 1635444444
transform 1 0 4324 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1635444444
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_29
timestamp 1635444444
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1635444444
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_47
timestamp 1635444444
transform 1 0 5428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_80_41
timestamp 1635444444
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1635444444
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1635444444
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_53
timestamp 1635444444
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1635444444
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1635444444
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_65
timestamp 1635444444
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1635444444
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1635444444
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1635444444
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1635444444
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1635444444
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_93
timestamp 1635444444
transform 1 0 9660 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_99
timestamp 1635444444
transform 1 0 10212 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_97
timestamp 1635444444
transform 1 0 10028 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1635444444
transform 1 0 9844 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1635444444
transform -1 0 10856 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1635444444
transform -1 0 10856 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_11
timestamp 1635444444
transform 1 0 2116 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1635444444
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1635444444
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _136_
timestamp 1635444444
transform -1 0 2484 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1635444444
transform -1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_15
timestamp 1635444444
transform 1 0 2484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_22
timestamp 1635444444
transform 1 0 3128 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _260_
timestamp 1635444444
transform -1 0 3128 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_34
timestamp 1635444444
transform 1 0 4232 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_46
timestamp 1635444444
transform 1 0 5336 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1635444444
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1635444444
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1635444444
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1635444444
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1635444444
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_93
timestamp 1635444444
transform 1 0 9660 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_99
timestamp 1635444444
transform 1 0 10212 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1635444444
transform 1 0 9844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1635444444
transform -1 0 10856 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_7
timestamp 1635444444
transform 1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1635444444
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _128_
timestamp 1635444444
transform 1 0 2116 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1635444444
transform -1 0 1748 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_14
timestamp 1635444444
transform 1 0 2392 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_22
timestamp 1635444444
transform 1 0 3128 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _168_
timestamp 1635444444
transform 1 0 2760 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_29
timestamp 1635444444
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1635444444
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_41
timestamp 1635444444
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_53
timestamp 1635444444
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_65
timestamp 1635444444
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1635444444
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1635444444
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_85
timestamp 1635444444
transform 1 0 8924 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1635444444
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_93
timestamp 1635444444
transform 1 0 9660 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_99
timestamp 1635444444
transform 1 0 10212 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1635444444
transform 1 0 9844 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1635444444
transform -1 0 10856 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_7
timestamp 1635444444
transform 1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1635444444
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1635444444
transform -1 0 1748 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1635444444
transform -1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_15
timestamp 1635444444
transform 1 0 2484 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_22
timestamp 1635444444
transform 1 0 3128 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _314_
timestamp 1635444444
transform 1 0 2852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_34
timestamp 1635444444
transform 1 0 4232 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_46
timestamp 1635444444
transform 1 0 5336 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_54
timestamp 1635444444
transform 1 0 6072 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_57
timestamp 1635444444
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1635444444
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_69
timestamp 1635444444
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_81
timestamp 1635444444
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_93
timestamp 1635444444
transform 1 0 9660 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_99
timestamp 1635444444
transform 1 0 10212 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1635444444
transform 1 0 9844 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1635444444
transform -1 0 10856 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_7
timestamp 1635444444
transform 1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1635444444
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _154_
timestamp 1635444444
transform -1 0 2392 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1635444444
transform -1 0 1748 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_14
timestamp 1635444444
transform 1 0 2392 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1635444444
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _259_
timestamp 1635444444
transform -1 0 3036 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1635444444
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_29
timestamp 1635444444
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1635444444
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_41
timestamp 1635444444
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_53
timestamp 1635444444
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_65
timestamp 1635444444
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1635444444
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1635444444
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_85
timestamp 1635444444
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1635444444
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_97
timestamp 1635444444
transform 1 0 10028 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1635444444
transform -1 0 10856 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_7
timestamp 1635444444
transform 1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_10
timestamp 1635444444
transform 1 0 2024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1635444444
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1635444444
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform -1 0 2024 0 1 48960
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1635444444
transform -1 0 1748 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1635444444
transform -1 0 2484 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_15
timestamp 1635444444
transform 1 0 2484 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_86_18
timestamp 1635444444
transform 1 0 2760 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1635444444
transform -1 0 3496 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1635444444
transform -1 0 2760 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_26
timestamp 1635444444
transform 1 0 3496 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_38
timestamp 1635444444
transform 1 0 4600 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_26
timestamp 1635444444
transform 1 0 3496 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_32
timestamp 1635444444
transform 1 0 4048 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1635444444
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _255_
timestamp 1635444444
transform -1 0 4048 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_85_50
timestamp 1635444444
transform 1 0 5704 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_86_44
timestamp 1635444444
transform 1 0 5152 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_57
timestamp 1635444444
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_56
timestamp 1635444444
transform 1 0 6256 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1635444444
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_69
timestamp 1635444444
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_68
timestamp 1635444444
transform 1 0 7360 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_81
timestamp 1635444444
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_80
timestamp 1635444444
transform 1 0 8464 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_85
timestamp 1635444444
transform 1 0 8924 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1635444444
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_93
timestamp 1635444444
transform 1 0 9660 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_99
timestamp 1635444444
transform 1 0 10212 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_93
timestamp 1635444444
transform 1 0 9660 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_99
timestamp 1635444444
transform 1 0 10212 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1635444444
transform 1 0 9844 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1635444444
transform 1 0 9844 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1635444444
transform -1 0 10856 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1635444444
transform -1 0 10856 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_87_10
timestamp 1635444444
transform 1 0 2024 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1635444444
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _172_
timestamp 1635444444
transform 1 0 1380 0 -1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_87_18
timestamp 1635444444
transform 1 0 2760 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _257_
timestamp 1635444444
transform -1 0 3588 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1635444444
transform 1 0 2392 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1635444444
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1635444444
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1635444444
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1635444444
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_57
timestamp 1635444444
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1635444444
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_69
timestamp 1635444444
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_81
timestamp 1635444444
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_101
timestamp 1635444444
transform 1 0 10396 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_87_93
timestamp 1635444444
transform 1 0 9660 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1635444444
transform -1 0 10856 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_88_10
timestamp 1635444444
transform 1 0 2024 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1635444444
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _175_
timestamp 1635444444
transform 1 0 1380 0 1 50048
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_88_24
timestamp 1635444444
transform 1 0 3312 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _138_
timestamp 1635444444
transform 1 0 2392 0 1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_88_32
timestamp 1635444444
transform 1 0 4048 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1635444444
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _256_
timestamp 1635444444
transform -1 0 4048 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _263_
timestamp 1635444444
transform -1 0 4692 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_39
timestamp 1635444444
transform 1 0 4692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_51
timestamp 1635444444
transform 1 0 5796 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_63
timestamp 1635444444
transform 1 0 6900 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_75
timestamp 1635444444
transform 1 0 8004 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1635444444
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_85
timestamp 1635444444
transform 1 0 8924 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1635444444
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_93
timestamp 1635444444
transform 1 0 9660 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_99
timestamp 1635444444
transform 1 0 10212 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1635444444
transform 1 0 9844 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1635444444
transform -1 0 10856 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_89_7
timestamp 1635444444
transform 1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1635444444
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 1635444444
transform 1 0 2116 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1635444444
transform -1 0 1748 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_14
timestamp 1635444444
transform 1 0 2392 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_21
timestamp 1635444444
transform 1 0 3036 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _141_
timestamp 1635444444
transform 1 0 2760 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _262_
timestamp 1635444444
transform -1 0 3680 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_28
timestamp 1635444444
transform 1 0 3680 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_40
timestamp 1635444444
transform 1 0 4784 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_52
timestamp 1635444444
transform 1 0 5888 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_57
timestamp 1635444444
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1635444444
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_69
timestamp 1635444444
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_81
timestamp 1635444444
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_93
timestamp 1635444444
transform 1 0 9660 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_99
timestamp 1635444444
transform 1 0 10212 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1635444444
transform 1 0 9844 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1635444444
transform -1 0 10856 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_7
timestamp 1635444444
transform 1 0 1748 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1635444444
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1635444444
transform -1 0 1748 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1635444444
transform -1 0 2484 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_90_15
timestamp 1635444444
transform 1 0 2484 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_22
timestamp 1635444444
transform 1 0 3128 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _147_
timestamp 1635444444
transform 1 0 2852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_29
timestamp 1635444444
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1635444444
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_41
timestamp 1635444444
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_53
timestamp 1635444444
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_65
timestamp 1635444444
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1635444444
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1635444444
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_85
timestamp 1635444444
transform 1 0 8924 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1635444444
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_93
timestamp 1635444444
transform 1 0 9660 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_99
timestamp 1635444444
transform 1 0 10212 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1635444444
transform 1 0 9844 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1635444444
transform -1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_7
timestamp 1635444444
transform 1 0 1748 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1635444444
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1635444444
transform -1 0 1748 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_91_22
timestamp 1635444444
transform 1 0 3128 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _264_
timestamp 1635444444
transform -1 0 3128 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_29
timestamp 1635444444
transform 1 0 3772 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _265_
timestamp 1635444444
transform -1 0 3772 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_41
timestamp 1635444444
transform 1 0 4876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1635444444
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_57
timestamp 1635444444
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1635444444
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_69
timestamp 1635444444
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_81
timestamp 1635444444
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_101
timestamp 1635444444
transform 1 0 10396 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_93
timestamp 1635444444
transform 1 0 9660 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1635444444
transform -1 0 10856 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_7
timestamp 1635444444
transform 1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_7
timestamp 1635444444
transform 1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1635444444
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1635444444
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _143_
timestamp 1635444444
transform 1 0 2116 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1635444444
transform -1 0 1748 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1635444444
transform -1 0 1748 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1635444444
transform -1 0 2484 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_92_14
timestamp 1635444444
transform 1 0 2392 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_92_21
timestamp 1635444444
transform 1 0 3036 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_93_15
timestamp 1635444444
transform 1 0 2484 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_93_23
timestamp 1635444444
transform 1 0 3220 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _266_
timestamp 1635444444
transform -1 0 3036 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1635444444
transform 1 0 2852 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1635444444
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_29
timestamp 1635444444
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_35
timestamp 1635444444
transform 1 0 4324 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1635444444
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_41
timestamp 1635444444
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1635444444
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_53
timestamp 1635444444
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1635444444
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_57
timestamp 1635444444
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1635444444
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_65
timestamp 1635444444
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1635444444
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_69
timestamp 1635444444
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1635444444
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_85
timestamp 1635444444
transform 1 0 8924 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_81
timestamp 1635444444
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1635444444
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_93
timestamp 1635444444
transform 1 0 9660 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_92_99
timestamp 1635444444
transform 1 0 10212 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_93
timestamp 1635444444
transform 1 0 9660 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_93_99
timestamp 1635444444
transform 1 0 10212 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1635444444
transform 1 0 9844 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1635444444
transform 1 0 9844 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1635444444
transform -1 0 10856 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1635444444
transform -1 0 10856 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_11
timestamp 1635444444
transform 1 0 2116 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1635444444
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1635444444
transform 1 0 1380 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_94_19
timestamp 1635444444
transform 1 0 2852 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1635444444
transform 1 0 2484 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1635444444
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_29
timestamp 1635444444
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1635444444
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_41
timestamp 1635444444
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_53
timestamp 1635444444
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_65
timestamp 1635444444
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1635444444
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1635444444
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_85
timestamp 1635444444
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1635444444
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_94_97
timestamp 1635444444
transform 1 0 10028 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1635444444
transform -1 0 10856 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_3
timestamp 1635444444
transform 1 0 1380 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1635444444
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _170_
timestamp 1635444444
transform 1 0 1564 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_95_15
timestamp 1635444444
transform 1 0 2484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_95_22
timestamp 1635444444
transform 1 0 3128 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _145_
timestamp 1635444444
transform 1 0 2852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_34
timestamp 1635444444
transform 1 0 4232 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_46
timestamp 1635444444
transform 1 0 5336 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1635444444
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_57
timestamp 1635444444
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1635444444
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_69
timestamp 1635444444
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_81
timestamp 1635444444
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_93
timestamp 1635444444
transform 1 0 9660 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_99
timestamp 1635444444
transform 1 0 10212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1635444444
transform 1 0 9844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1635444444
transform -1 0 10856 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_7
timestamp 1635444444
transform 1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1635444444
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1635444444
transform -1 0 1748 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1635444444
transform -1 0 2484 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1635444444
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1635444444
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_29
timestamp 1635444444
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1635444444
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_41
timestamp 1635444444
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_53
timestamp 1635444444
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_65
timestamp 1635444444
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1635444444
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1635444444
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_85
timestamp 1635444444
transform 1 0 8924 0 1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1635444444
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_93
timestamp 1635444444
transform 1 0 9660 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_96_99
timestamp 1635444444
transform 1 0 10212 0 1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1635444444
transform 1 0 9936 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1635444444
transform -1 0 10856 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_11
timestamp 1635444444
transform 1 0 2116 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1635444444
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _174_
timestamp 1635444444
transform 1 0 1380 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_97_19
timestamp 1635444444
transform 1 0 2852 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1635444444
transform 1 0 2484 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_97_31
timestamp 1635444444
transform 1 0 3956 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_43
timestamp 1635444444
transform 1 0 5060 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1635444444
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_57
timestamp 1635444444
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1635444444
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_69
timestamp 1635444444
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_81
timestamp 1635444444
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_97_93
timestamp 1635444444
transform 1 0 9660 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_97_99
timestamp 1635444444
transform 1 0 10212 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1635444444
transform 1 0 9936 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1635444444
transform -1 0 10856 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_98_11
timestamp 1635444444
transform 1 0 2116 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_7
timestamp 1635444444
transform 1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1635444444
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _169_
timestamp 1635444444
transform 1 0 2208 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1635444444
transform -1 0 1748 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_16
timestamp 1635444444
transform 1 0 2576 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_24
timestamp 1635444444
transform 1 0 3312 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1635444444
transform 1 0 2944 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_33
timestamp 1635444444
transform 1 0 4140 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1635444444
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1635444444
transform 1 0 3772 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_45
timestamp 1635444444
transform 1 0 5244 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_57
timestamp 1635444444
transform 1 0 6348 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_69
timestamp 1635444444
transform 1 0 7452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_81
timestamp 1635444444
transform 1 0 8556 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_85
timestamp 1635444444
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1635444444
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_97
timestamp 1635444444
transform 1 0 10028 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1635444444
transform -1 0 10856 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_100_7
timestamp 1635444444
transform 1 0 1748 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_11
timestamp 1635444444
transform 1 0 2116 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_7
timestamp 1635444444
transform 1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1635444444
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1635444444
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1635444444
transform -1 0 2576 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1635444444
transform -1 0 1748 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1635444444
transform -1 0 1748 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_20
timestamp 1635444444
transform 1 0 2944 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_16
timestamp 1635444444
transform 1 0 2576 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_24
timestamp 1635444444
transform 1 0 3312 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _189_
timestamp 1635444444
transform 1 0 2300 0 1 56576
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1635444444
transform 1 0 2944 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_29
timestamp 1635444444
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_36
timestamp 1635444444
transform 1 0 4416 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1635444444
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_41
timestamp 1635444444
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_48
timestamp 1635444444
transform 1 0 5520 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_53
timestamp 1635444444
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_57
timestamp 1635444444
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1635444444
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_65
timestamp 1635444444
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1635444444
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_99_69
timestamp 1635444444
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1635444444
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_100_85
timestamp 1635444444
transform 1 0 8924 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_81
timestamp 1635444444
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1635444444
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1635444444
transform -1 0 10212 0 1 56576
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_100_99
timestamp 1635444444
transform 1 0 10212 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_99_93
timestamp 1635444444
transform 1 0 9660 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_99
timestamp 1635444444
transform 1 0 10212 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1635444444
transform 1 0 9936 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1635444444
transform -1 0 10856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1635444444
transform -1 0 10856 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_11
timestamp 1635444444
transform 1 0 2116 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1635444444
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _179_
timestamp 1635444444
transform 1 0 1380 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_101_22
timestamp 1635444444
transform 1 0 3128 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _188_
timestamp 1635444444
transform -1 0 3128 0 -1 57664
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_101_34
timestamp 1635444444
transform 1 0 4232 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_46
timestamp 1635444444
transform 1 0 5336 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1635444444
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_57
timestamp 1635444444
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1635444444
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_69
timestamp 1635444444
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_81
timestamp 1635444444
transform 1 0 8556 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_101
timestamp 1635444444
transform 1 0 10396 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_93
timestamp 1635444444
transform 1 0 9660 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1635444444
transform -1 0 10856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_11
timestamp 1635444444
transform 1 0 2116 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1635444444
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _178_
timestamp 1635444444
transform 1 0 1380 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_102_19
timestamp 1635444444
transform 1 0 2852 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1635444444
transform -1 0 2852 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 1635444444
transform 1 0 3588 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_29
timestamp 1635444444
transform 1 0 3772 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1635444444
transform 1 0 3680 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_41
timestamp 1635444444
transform 1 0 4876 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_53
timestamp 1635444444
transform 1 0 5980 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_65
timestamp 1635444444
transform 1 0 7084 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_102_77
timestamp 1635444444
transform 1 0 8188 0 1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_102_83
timestamp 1635444444
transform 1 0 8740 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_85
timestamp 1635444444
transform 1 0 8924 0 1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1635444444
transform 1 0 8832 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_102_93
timestamp 1635444444
transform 1 0 9660 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_102_99
timestamp 1635444444
transform 1 0 10212 0 1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1635444444
transform 1 0 9936 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1635444444
transform -1 0 10856 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_103_7
timestamp 1635444444
transform 1 0 1748 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1635444444
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1635444444
transform -1 0 1748 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_103_19
timestamp 1635444444
transform 1 0 2852 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_31
timestamp 1635444444
transform 1 0 3956 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_43
timestamp 1635444444
transform 1 0 5060 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_55
timestamp 1635444444
transform 1 0 6164 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_57
timestamp 1635444444
transform 1 0 6348 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1635444444
transform 1 0 6256 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_69
timestamp 1635444444
transform 1 0 7452 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_81
timestamp 1635444444
transform 1 0 8556 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_103_93
timestamp 1635444444
transform 1 0 9660 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_103_99
timestamp 1635444444
transform 1 0 10212 0 -1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1635444444
transform 1 0 9936 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1635444444
transform -1 0 10856 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_7
timestamp 1635444444
transform 1 0 1748 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1635444444
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _177_
timestamp 1635444444
transform 1 0 2116 0 1 58752
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1635444444
transform -1 0 1748 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_104_21
timestamp 1635444444
transform 1 0 3036 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 1635444444
transform 1 0 3588 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_29
timestamp 1635444444
transform 1 0 3772 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1635444444
transform 1 0 3680 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_41
timestamp 1635444444
transform 1 0 4876 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_53
timestamp 1635444444
transform 1 0 5980 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_65
timestamp 1635444444
transform 1 0 7084 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_104_77
timestamp 1635444444
transform 1 0 8188 0 1 58752
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_83
timestamp 1635444444
transform 1 0 8740 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_85
timestamp 1635444444
transform 1 0 8924 0 1 58752
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1635444444
transform 1 0 8832 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_93
timestamp 1635444444
transform 1 0 9660 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_104_99
timestamp 1635444444
transform 1 0 10212 0 1 58752
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1635444444
transform 1 0 9936 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1635444444
transform -1 0 10856 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_105_7
timestamp 1635444444
transform 1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_11
timestamp 1635444444
transform 1 0 2116 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_106_7
timestamp 1635444444
transform 1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1635444444
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1635444444
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _176_
timestamp 1635444444
transform 1 0 2208 0 1 59840
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1635444444
transform -1 0 1748 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1635444444
transform -1 0 1748 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1635444444
transform 1 0 2116 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1635444444
transform 1 0 2484 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_22
timestamp 1635444444
transform 1 0 3128 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1635444444
transform 1 0 3588 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_29
timestamp 1635444444
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1635444444
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1635444444
transform 1 0 4692 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_51
timestamp 1635444444
transform 1 0 5796 0 -1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_41
timestamp 1635444444
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_55
timestamp 1635444444
transform 1 0 6164 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_57
timestamp 1635444444
transform 1 0 6348 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_53
timestamp 1635444444
transform 1 0 5980 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1635444444
transform 1 0 6256 0 -1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_69
timestamp 1635444444
transform 1 0 7452 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_65
timestamp 1635444444
transform 1 0 7084 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_77
timestamp 1635444444
transform 1 0 8188 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_105_81
timestamp 1635444444
transform 1 0 8556 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_83
timestamp 1635444444
transform 1 0 8740 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_85
timestamp 1635444444
transform 1 0 8924 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1635444444
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_105_101
timestamp 1635444444
transform 1 0 10396 0 -1 59840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_105_93
timestamp 1635444444
transform 1 0 9660 0 -1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_93
timestamp 1635444444
transform 1 0 9660 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_106_99
timestamp 1635444444
transform 1 0 10212 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1635444444
transform 1 0 9936 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1635444444
transform -1 0 10856 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1635444444
transform -1 0 10856 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_107_7
timestamp 1635444444
transform 1 0 1748 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1635444444
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1635444444
transform -1 0 1748 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_107_21
timestamp 1635444444
transform 1 0 3036 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_2  _185_
timestamp 1635444444
transform 1 0 2300 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_107_33
timestamp 1635444444
transform 1 0 4140 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_45
timestamp 1635444444
transform 1 0 5244 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_53
timestamp 1635444444
transform 1 0 5980 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_57
timestamp 1635444444
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1635444444
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_69
timestamp 1635444444
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_81
timestamp 1635444444
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_93
timestamp 1635444444
transform 1 0 9660 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_107_99
timestamp 1635444444
transform 1 0 10212 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1635444444
transform 1 0 9936 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1635444444
transform -1 0 10856 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_108_11
timestamp 1635444444
transform 1 0 2116 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1635444444
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 1635444444
transform -1 0 2116 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_108_19
timestamp 1635444444
transform 1 0 2852 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1635444444
transform 1 0 2484 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1635444444
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_33
timestamp 1635444444
transform 1 0 4140 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1635444444
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1635444444
transform 1 0 3772 0 1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_45
timestamp 1635444444
transform 1 0 5244 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_57
timestamp 1635444444
transform 1 0 6348 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_69
timestamp 1635444444
transform 1 0 7452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_108_81
timestamp 1635444444
transform 1 0 8556 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_85
timestamp 1635444444
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1635444444
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_108_97
timestamp 1635444444
transform 1 0 10028 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1635444444
transform -1 0 10856 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_11
timestamp 1635444444
transform 1 0 2116 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1635444444
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _182_
timestamp 1635444444
transform 1 0 1380 0 -1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_109_19
timestamp 1635444444
transform 1 0 2852 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1635444444
transform 1 0 2484 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_109_31
timestamp 1635444444
transform 1 0 3956 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_43
timestamp 1635444444
transform 1 0 5060 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1635444444
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_57
timestamp 1635444444
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1635444444
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_69
timestamp 1635444444
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_81
timestamp 1635444444
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_109_93
timestamp 1635444444
transform 1 0 9660 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_109_99
timestamp 1635444444
transform 1 0 10212 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1635444444
transform 1 0 9936 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1635444444
transform -1 0 10856 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_11
timestamp 1635444444
transform 1 0 2116 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1635444444
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _181_
timestamp 1635444444
transform 1 0 1380 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_110_23
timestamp 1635444444
transform 1 0 3220 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 1635444444
transform -1 0 3220 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1635444444
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_29
timestamp 1635444444
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1635444444
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_41
timestamp 1635444444
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_53
timestamp 1635444444
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_65
timestamp 1635444444
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1635444444
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1635444444
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_85
timestamp 1635444444
transform 1 0 8924 0 1 62016
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1635444444
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_110_93
timestamp 1635444444
transform 1 0 9660 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_110_99
timestamp 1635444444
transform 1 0 10212 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1635444444
transform 1 0 9936 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1635444444
transform -1 0 10856 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_7
timestamp 1635444444
transform 1 0 1748 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1635444444
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1635444444
transform -1 0 1748 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1635444444
transform -1 0 2484 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_111_15
timestamp 1635444444
transform 1 0 2484 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _183_
timestamp 1635444444
transform 1 0 2852 0 -1 63104
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_111_29
timestamp 1635444444
transform 1 0 3772 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_36
timestamp 1635444444
transform 1 0 4416 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 1635444444
transform 1 0 4140 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_111_48
timestamp 1635444444
transform 1 0 5520 0 -1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_111_57
timestamp 1635444444
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1635444444
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_69
timestamp 1635444444
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_81
timestamp 1635444444
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_93
timestamp 1635444444
transform 1 0 9660 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_111_99
timestamp 1635444444
transform 1 0 10212 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1635444444
transform 1 0 9936 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1635444444
transform -1 0 10856 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_112_11
timestamp 1635444444
transform 1 0 2116 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_3
timestamp 1635444444
transform 1 0 1380 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_7
timestamp 1635444444
transform 1 0 1748 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1635444444
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1635444444
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _192_
timestamp 1635444444
transform 1 0 1380 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _193_
timestamp 1635444444
transform -1 0 2576 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_112_23
timestamp 1635444444
transform 1 0 3220 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_16
timestamp 1635444444
transform 1 0 2576 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_113_24
timestamp 1635444444
transform 1 0 3312 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _187_
timestamp 1635444444
transform -1 0 3220 0 1 63104
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1635444444
transform 1 0 2944 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1635444444
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_33
timestamp 1635444444
transform 1 0 4140 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_32
timestamp 1635444444
transform 1 0 4048 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1635444444
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1635444444
transform 1 0 3772 0 1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1635444444
transform 1 0 3680 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_112_45
timestamp 1635444444
transform 1 0 5244 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_44
timestamp 1635444444
transform 1 0 5152 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_57
timestamp 1635444444
transform 1 0 6348 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_57
timestamp 1635444444
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1635444444
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_69
timestamp 1635444444
transform 1 0 7452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_69
timestamp 1635444444
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_112_81
timestamp 1635444444
transform 1 0 8556 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_85
timestamp 1635444444
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_81
timestamp 1635444444
transform 1 0 8556 0 -1 64192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1635444444
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1635444444
transform -1 0 10212 0 -1 64192
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_112_97
timestamp 1635444444
transform 1 0 10028 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_113_99
timestamp 1635444444
transform 1 0 10212 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1635444444
transform -1 0 10856 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1635444444
transform -1 0 10856 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_114_7
timestamp 1635444444
transform 1 0 1748 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1635444444
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1635444444
transform -1 0 1748 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_114_23
timestamp 1635444444
transform 1 0 3220 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _191_
timestamp 1635444444
transform 1 0 2300 0 1 64192
box -38 -48 958 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1635444444
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_29
timestamp 1635444444
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1635444444
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_41
timestamp 1635444444
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_53
timestamp 1635444444
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_65
timestamp 1635444444
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1635444444
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1635444444
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_114_85
timestamp 1635444444
transform 1 0 8924 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1635444444
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1635444444
transform -1 0 10212 0 1 64192
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_114_99
timestamp 1635444444
transform 1 0 10212 0 1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1635444444
transform -1 0 10856 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_115_3
timestamp 1635444444
transform 1 0 1380 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1635444444
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _194_
timestamp 1635444444
transform 1 0 1748 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_115_15
timestamp 1635444444
transform 1 0 2484 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _190_
timestamp 1635444444
transform 1 0 2852 0 -1 65280
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_115_29
timestamp 1635444444
transform 1 0 3772 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_41
timestamp 1635444444
transform 1 0 4876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_115_53
timestamp 1635444444
transform 1 0 5980 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_57
timestamp 1635444444
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1635444444
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_69
timestamp 1635444444
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_81
timestamp 1635444444
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_115_101
timestamp 1635444444
transform 1 0 10396 0 -1 65280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_115_93
timestamp 1635444444
transform 1 0 9660 0 -1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1635444444
transform -1 0 10856 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_7
timestamp 1635444444
transform 1 0 1748 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1635444444
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1635444444
transform -1 0 1748 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1635444444
transform 1 0 2116 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_15
timestamp 1635444444
transform 1 0 2484 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_116_23
timestamp 1635444444
transform 1 0 3220 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1635444444
transform 1 0 2852 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1635444444
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_29
timestamp 1635444444
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1635444444
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_41
timestamp 1635444444
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_53
timestamp 1635444444
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_65
timestamp 1635444444
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1635444444
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1635444444
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_85
timestamp 1635444444
transform 1 0 8924 0 1 65280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1635444444
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_116_93
timestamp 1635444444
transform 1 0 9660 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_116_99
timestamp 1635444444
transform 1 0 10212 0 1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1635444444
transform 1 0 9936 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1635444444
transform -1 0 10856 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1635444444
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1635444444
transform 1 0 1380 0 -1 66368
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_117_13
timestamp 1635444444
transform 1 0 2300 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_25
timestamp 1635444444
transform 1 0 3404 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_37
timestamp 1635444444
transform 1 0 4508 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_49
timestamp 1635444444
transform 1 0 5612 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1635444444
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_57
timestamp 1635444444
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1635444444
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_69
timestamp 1635444444
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_81
timestamp 1635444444
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_117_93
timestamp 1635444444
transform 1 0 9660 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_117_99
timestamp 1635444444
transform 1 0 10212 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1635444444
transform 1 0 9936 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1635444444
transform -1 0 10856 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_7
timestamp 1635444444
transform 1 0 1748 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_119_3
timestamp 1635444444
transform 1 0 1380 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1635444444
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1635444444
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _195_
timestamp 1635444444
transform -1 0 2484 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1635444444
transform 1 0 2116 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1635444444
transform -1 0 1748 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_118_14
timestamp 1635444444
transform 1 0 2392 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_118_21
timestamp 1635444444
transform 1 0 3036 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_119_15
timestamp 1635444444
transform 1 0 2484 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_119_23
timestamp 1635444444
transform 1 0 3220 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _197_
timestamp 1635444444
transform -1 0 3220 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1635444444
transform 1 0 2760 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1635444444
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_29
timestamp 1635444444
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_35
timestamp 1635444444
transform 1 0 4324 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1635444444
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_41
timestamp 1635444444
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_47
timestamp 1635444444
transform 1 0 5428 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_118_53
timestamp 1635444444
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1635444444
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_57
timestamp 1635444444
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1635444444
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_65
timestamp 1635444444
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1635444444
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_119_69
timestamp 1635444444
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1635444444
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_85
timestamp 1635444444
transform 1 0 8924 0 1 66368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_119_81
timestamp 1635444444
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1635444444
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_118_93
timestamp 1635444444
transform 1 0 9660 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_118_99
timestamp 1635444444
transform 1 0 10212 0 1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_119_101
timestamp 1635444444
transform 1 0 10396 0 -1 67456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_119_93
timestamp 1635444444
transform 1 0 9660 0 -1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1635444444
transform 1 0 9936 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1635444444
transform -1 0 10856 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1635444444
transform -1 0 10856 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1635444444
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1635444444
transform 1 0 1380 0 1 67456
box -38 -48 958 592
use sky130_fd_sc_hd__decap_6  FILLER_120_13
timestamp 1635444444
transform 1 0 2300 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_120_23
timestamp 1635444444
transform 1 0 3220 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1635444444
transform 1 0 2852 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1635444444
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_29
timestamp 1635444444
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1635444444
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_41
timestamp 1635444444
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_53
timestamp 1635444444
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_65
timestamp 1635444444
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1635444444
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1635444444
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_85
timestamp 1635444444
transform 1 0 8924 0 1 67456
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1635444444
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_120_93
timestamp 1635444444
transform 1 0 9660 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_120_99
timestamp 1635444444
transform 1 0 10212 0 1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1635444444
transform 1 0 9936 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1635444444
transform -1 0 10856 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_3
timestamp 1635444444
transform 1 0 1380 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1635444444
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _196_
timestamp 1635444444
transform 1 0 1748 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_121_15
timestamp 1635444444
transform 1 0 2484 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _199_
timestamp 1635444444
transform 1 0 2852 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_121_27
timestamp 1635444444
transform 1 0 3588 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_121_34
timestamp 1635444444
transform 1 0 4232 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1635444444
transform 1 0 3956 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_121_46
timestamp 1635444444
transform 1 0 5336 0 -1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_54
timestamp 1635444444
transform 1 0 6072 0 -1 68544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_57
timestamp 1635444444
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1635444444
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_69
timestamp 1635444444
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_81
timestamp 1635444444
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_93
timestamp 1635444444
transform 1 0 9660 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_121_99
timestamp 1635444444
transform 1 0 10212 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1635444444
transform 1 0 9936 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1635444444
transform -1 0 10856 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_6
timestamp 1635444444
transform 1 0 1656 0 1 68544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1635444444
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1635444444
transform -1 0 1656 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_122_24
timestamp 1635444444
transform 1 0 3312 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _204_
timestamp 1635444444
transform -1 0 3312 0 1 68544
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_122_32
timestamp 1635444444
transform 1 0 4048 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1635444444
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1635444444
transform 1 0 3772 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_44
timestamp 1635444444
transform 1 0 5152 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_56
timestamp 1635444444
transform 1 0 6256 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_68
timestamp 1635444444
transform 1 0 7360 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_122_80
timestamp 1635444444
transform 1 0 8464 0 1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_85
timestamp 1635444444
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1635444444
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_122_97
timestamp 1635444444
transform 1 0 10028 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1635444444
transform -1 0 10856 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_123_11
timestamp 1635444444
transform 1 0 2116 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1635444444
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _200_
timestamp 1635444444
transform -1 0 2116 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_17
timestamp 1635444444
transform 1 0 2668 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _205_
timestamp 1635444444
transform 1 0 2760 0 -1 69632
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_123_28
timestamp 1635444444
transform 1 0 3680 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_35
timestamp 1635444444
transform 1 0 4324 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1635444444
transform 1 0 4048 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_123_47
timestamp 1635444444
transform 1 0 5428 0 -1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1635444444
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_57
timestamp 1635444444
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1635444444
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_69
timestamp 1635444444
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_81
timestamp 1635444444
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_93
timestamp 1635444444
transform 1 0 9660 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_123_99
timestamp 1635444444
transform 1 0 10212 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1635444444
transform 1 0 9936 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1635444444
transform -1 0 10856 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_124_12
timestamp 1635444444
transform 1 0 2208 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_124_6
timestamp 1635444444
transform 1 0 1656 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1635444444
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1635444444
transform -1 0 1656 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_124_21
timestamp 1635444444
transform 1 0 3036 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _206_
timestamp 1635444444
transform -1 0 3036 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1635444444
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_32
timestamp 1635444444
transform 1 0 4048 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1635444444
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1635444444
transform 1 0 3772 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_44
timestamp 1635444444
transform 1 0 5152 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_56
timestamp 1635444444
transform 1 0 6256 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_68
timestamp 1635444444
transform 1 0 7360 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_124_80
timestamp 1635444444
transform 1 0 8464 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_124_85
timestamp 1635444444
transform 1 0 8924 0 1 69632
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1635444444
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_124_93
timestamp 1635444444
transform 1 0 9660 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_124_99
timestamp 1635444444
transform 1 0 10212 0 1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1635444444
transform 1 0 9936 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1635444444
transform -1 0 10856 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_125_3
timestamp 1635444444
transform 1 0 1380 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_125_8
timestamp 1635444444
transform 1 0 1840 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1635444444
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1635444444
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1635444444
transform -1 0 1840 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _207_
timestamp 1635444444
transform -1 0 2944 0 -1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1635444444
transform 1 0 1380 0 1 70720
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_125_20
timestamp 1635444444
transform 1 0 2944 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_126_13
timestamp 1635444444
transform 1 0 2300 0 1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_126_20
timestamp 1635444444
transform 1 0 2944 0 1 70720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1635444444
transform -1 0 2944 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1635444444
transform 1 0 3312 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_27
timestamp 1635444444
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_29
timestamp 1635444444
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1635444444
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_39
timestamp 1635444444
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1635444444
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_41
timestamp 1635444444
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1635444444
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_57
timestamp 1635444444
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_53
timestamp 1635444444
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1635444444
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_69
timestamp 1635444444
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_65
timestamp 1635444444
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1635444444
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_125_81
timestamp 1635444444
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1635444444
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_126_85
timestamp 1635444444
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1635444444
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_125_93
timestamp 1635444444
transform 1 0 9660 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_125_99
timestamp 1635444444
transform 1 0 10212 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_126_97
timestamp 1635444444
transform 1 0 10028 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1635444444
transform 1 0 9936 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1635444444
transform -1 0 10856 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1635444444
transform -1 0 10856 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1635444444
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1635444444
transform 1 0 1380 0 -1 71808
box -38 -48 958 592
use sky130_fd_sc_hd__decap_12  FILLER_127_13
timestamp 1635444444
transform 1 0 2300 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_25
timestamp 1635444444
transform 1 0 3404 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_37
timestamp 1635444444
transform 1 0 4508 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_49
timestamp 1635444444
transform 1 0 5612 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1635444444
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_57
timestamp 1635444444
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1635444444
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_69
timestamp 1635444444
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_81
timestamp 1635444444
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_127_93
timestamp 1635444444
transform 1 0 9660 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_127_99
timestamp 1635444444
transform 1 0 10212 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1635444444
transform 1 0 9936 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1635444444
transform -1 0 10856 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_11
timestamp 1635444444
transform 1 0 2116 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1635444444
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _201_
timestamp 1635444444
transform 1 0 1380 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_128_23
timestamp 1635444444
transform 1 0 3220 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1635444444
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_29
timestamp 1635444444
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1635444444
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_41
timestamp 1635444444
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_53
timestamp 1635444444
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_65
timestamp 1635444444
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1635444444
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1635444444
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_85
timestamp 1635444444
transform 1 0 8924 0 1 71808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1635444444
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_128_93
timestamp 1635444444
transform 1 0 9660 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_128_99
timestamp 1635444444
transform 1 0 10212 0 1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1635444444
transform 1 0 9936 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1635444444
transform -1 0 10856 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_6
timestamp 1635444444
transform 1 0 1656 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1635444444
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1635444444
transform -1 0 1656 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_18
timestamp 1635444444
transform 1 0 2760 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_30
timestamp 1635444444
transform 1 0 3864 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_42
timestamp 1635444444
transform 1 0 4968 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_54
timestamp 1635444444
transform 1 0 6072 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_57
timestamp 1635444444
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1635444444
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_69
timestamp 1635444444
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_81
timestamp 1635444444
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_101
timestamp 1635444444
transform 1 0 10396 0 -1 72896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_129_93
timestamp 1635444444
transform 1 0 9660 0 -1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1635444444
transform -1 0 10856 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_6
timestamp 1635444444
transform 1 0 1656 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1635444444
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1635444444
transform -1 0 1656 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1635444444
transform 1 0 2024 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_13
timestamp 1635444444
transform 1 0 2300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_130_25
timestamp 1635444444
transform 1 0 3404 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_29
timestamp 1635444444
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1635444444
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_41
timestamp 1635444444
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_53
timestamp 1635444444
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_65
timestamp 1635444444
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1635444444
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1635444444
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_85
timestamp 1635444444
transform 1 0 8924 0 1 72896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1635444444
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_130_93
timestamp 1635444444
transform 1 0 9660 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_130_99
timestamp 1635444444
transform 1 0 10212 0 1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1635444444
transform 1 0 9936 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1635444444
transform -1 0 10856 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_11
timestamp 1635444444
transform 1 0 2116 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1635444444
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _203_
timestamp 1635444444
transform -1 0 2116 0 -1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_131_18
timestamp 1635444444
transform 1 0 2760 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1635444444
transform 1 0 2484 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_30
timestamp 1635444444
transform 1 0 3864 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_42
timestamp 1635444444
transform 1 0 4968 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_54
timestamp 1635444444
transform 1 0 6072 0 -1 73984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_57
timestamp 1635444444
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1635444444
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_69
timestamp 1635444444
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_81
timestamp 1635444444
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_93
timestamp 1635444444
transform 1 0 9660 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_131_99
timestamp 1635444444
transform 1 0 10212 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1635444444
transform 1 0 9936 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1635444444
transform -1 0 10856 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_11
timestamp 1635444444
transform 1 0 2116 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_12
timestamp 1635444444
transform 1 0 2208 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_133_6
timestamp 1635444444
transform 1 0 1656 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1635444444
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1635444444
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _202_
timestamp 1635444444
transform 1 0 1380 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1635444444
transform -1 0 1656 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_23
timestamp 1635444444
transform 1 0 3220 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_133_21
timestamp 1635444444
transform 1 0 3036 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _208_
timestamp 1635444444
transform -1 0 3220 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _210_
timestamp 1635444444
transform -1 0 3036 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _211_
timestamp 1635444444
transform 1 0 3404 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1635444444
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_29
timestamp 1635444444
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_33
timestamp 1635444444
transform 1 0 4140 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1635444444
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_41
timestamp 1635444444
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_45
timestamp 1635444444
transform 1 0 5244 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_132_53
timestamp 1635444444
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_53
timestamp 1635444444
transform 1 0 5980 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_133_57
timestamp 1635444444
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1635444444
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_65
timestamp 1635444444
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1635444444
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_133_69
timestamp 1635444444
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1635444444
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_85
timestamp 1635444444
transform 1 0 8924 0 1 73984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_133_81
timestamp 1635444444
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1635444444
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_132_93
timestamp 1635444444
transform 1 0 9660 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_132_99
timestamp 1635444444
transform 1 0 10212 0 1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_133_101
timestamp 1635444444
transform 1 0 10396 0 -1 75072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_133_93
timestamp 1635444444
transform 1 0 9660 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1635444444
transform 1 0 9936 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1635444444
transform -1 0 10856 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1635444444
transform -1 0 10856 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_134_12
timestamp 1635444444
transform 1 0 2208 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_6
timestamp 1635444444
transform 1 0 1656 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1635444444
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1635444444
transform -1 0 1656 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_134_21
timestamp 1635444444
transform 1 0 3036 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _209_
timestamp 1635444444
transform -1 0 3036 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1635444444
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_32
timestamp 1635444444
transform 1 0 4048 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1635444444
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1635444444
transform 1 0 3772 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_44
timestamp 1635444444
transform 1 0 5152 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_56
timestamp 1635444444
transform 1 0 6256 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_68
timestamp 1635444444
transform 1 0 7360 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_134_80
timestamp 1635444444
transform 1 0 8464 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_134_85
timestamp 1635444444
transform 1 0 8924 0 1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1635444444
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_134_93
timestamp 1635444444
transform 1 0 9660 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_134_99
timestamp 1635444444
transform 1 0 10212 0 1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1635444444
transform 1 0 9936 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1635444444
transform -1 0 10856 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_135_3
timestamp 1635444444
transform 1 0 1380 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1635444444
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _212_
timestamp 1635444444
transform 1 0 1656 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_135_14
timestamp 1635444444
transform 1 0 2392 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_21
timestamp 1635444444
transform 1 0 3036 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1635444444
transform 1 0 2760 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_33
timestamp 1635444444
transform 1 0 4140 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_45
timestamp 1635444444
transform 1 0 5244 0 -1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_53
timestamp 1635444444
transform 1 0 5980 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_57
timestamp 1635444444
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1635444444
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_69
timestamp 1635444444
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_81
timestamp 1635444444
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_135_93
timestamp 1635444444
transform 1 0 9660 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_135_99
timestamp 1635444444
transform 1 0 10212 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1635444444
transform 1 0 9936 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1635444444
transform -1 0 10856 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_136_3
timestamp 1635444444
transform 1 0 1380 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1635444444
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _213_
timestamp 1635444444
transform 1 0 1656 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_136_14
timestamp 1635444444
transform 1 0 2392 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_136_21
timestamp 1635444444
transform 1 0 3036 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1635444444
transform 1 0 2760 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1635444444
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_29
timestamp 1635444444
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1635444444
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_41
timestamp 1635444444
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_53
timestamp 1635444444
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_65
timestamp 1635444444
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1635444444
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1635444444
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_85
timestamp 1635444444
transform 1 0 8924 0 1 76160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1635444444
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_136_93
timestamp 1635444444
transform 1 0 9660 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_136_99
timestamp 1635444444
transform 1 0 10212 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1635444444
transform 1 0 9936 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1635444444
transform -1 0 10856 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_6
timestamp 1635444444
transform 1 0 1656 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1635444444
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1635444444
transform -1 0 1656 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1635444444
transform -1 0 2300 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_13
timestamp 1635444444
transform 1 0 2300 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_137_20
timestamp 1635444444
transform 1 0 2944 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1635444444
transform -1 0 2944 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1635444444
transform -1 0 3588 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_27
timestamp 1635444444
transform 1 0 3588 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_137_34
timestamp 1635444444
transform 1 0 4232 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1635444444
transform 1 0 3956 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_137_46
timestamp 1635444444
transform 1 0 5336 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_137_54
timestamp 1635444444
transform 1 0 6072 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_137_57
timestamp 1635444444
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1635444444
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_69
timestamp 1635444444
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_81
timestamp 1635444444
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_93
timestamp 1635444444
transform 1 0 9660 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_137_99
timestamp 1635444444
transform 1 0 10212 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1635444444
transform 1 0 9936 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1635444444
transform -1 0 10856 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_11
timestamp 1635444444
transform 1 0 2116 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_3
timestamp 1635444444
transform 1 0 1380 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1635444444
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1635444444
transform -1 0 2116 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_18
timestamp 1635444444
transform 1 0 2760 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1635444444
transform -1 0 2760 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_138_26
timestamp 1635444444
transform 1 0 3496 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_138_32
timestamp 1635444444
transform 1 0 4048 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1635444444
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1635444444
transform 1 0 3772 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1635444444
transform 1 0 4416 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_39
timestamp 1635444444
transform 1 0 4692 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_138_46
timestamp 1635444444
transform 1 0 5336 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1635444444
transform 1 0 5060 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_138_54
timestamp 1635444444
transform 1 0 6072 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_138_57
timestamp 1635444444
transform 1 0 6348 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1635444444
transform 1 0 6256 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_69
timestamp 1635444444
transform 1 0 7452 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_138_81
timestamp 1635444444
transform 1 0 8556 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_138_85
timestamp 1635444444
transform 1 0 8924 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1635444444
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1635444444
transform 1 0 9200 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_138_91
timestamp 1635444444
transform 1 0 9476 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_138_99
timestamp 1635444444
transform 1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1635444444
transform -1 0 10212 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1635444444
transform -1 0 10856 0 1 77248
box -38 -48 314 592
<< labels >>
rlabel metal4 s 2575 2128 2895 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 5839 2128 6159 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 9103 2128 9423 77840 6 vccd1
port 0 nsew power input
rlabel metal4 s 4207 2128 4527 77840 6 vssd1
port 1 nsew ground input
rlabel metal4 s 7471 2128 7791 77840 6 vssd1
port 1 nsew ground input
rlabel metal3 s 11200 79432 12000 79552 6 wb_clk_i
port 2 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wb_rst_i
port 3 nsew signal input
rlabel metal3 s 11200 78616 12000 78736 6 wbm_a_ack_i
port 4 nsew signal input
rlabel metal3 s 11200 5584 12000 5704 6 wbm_a_adr_o[0]
port 5 nsew signal tristate
rlabel metal3 s 11200 13200 12000 13320 6 wbm_a_adr_o[10]
port 6 nsew signal tristate
rlabel metal3 s 11200 13880 12000 14000 6 wbm_a_adr_o[11]
port 7 nsew signal tristate
rlabel metal3 s 11200 14696 12000 14816 6 wbm_a_adr_o[12]
port 8 nsew signal tristate
rlabel metal3 s 11200 15512 12000 15632 6 wbm_a_adr_o[13]
port 9 nsew signal tristate
rlabel metal3 s 11200 16192 12000 16312 6 wbm_a_adr_o[14]
port 10 nsew signal tristate
rlabel metal3 s 11200 17008 12000 17128 6 wbm_a_adr_o[15]
port 11 nsew signal tristate
rlabel metal3 s 11200 17688 12000 17808 6 wbm_a_adr_o[16]
port 12 nsew signal tristate
rlabel metal3 s 11200 18504 12000 18624 6 wbm_a_adr_o[17]
port 13 nsew signal tristate
rlabel metal3 s 11200 19320 12000 19440 6 wbm_a_adr_o[18]
port 14 nsew signal tristate
rlabel metal3 s 11200 20000 12000 20120 6 wbm_a_adr_o[19]
port 15 nsew signal tristate
rlabel metal3 s 11200 6264 12000 6384 6 wbm_a_adr_o[1]
port 16 nsew signal tristate
rlabel metal3 s 11200 20816 12000 20936 6 wbm_a_adr_o[20]
port 17 nsew signal tristate
rlabel metal3 s 11200 21496 12000 21616 6 wbm_a_adr_o[21]
port 18 nsew signal tristate
rlabel metal3 s 11200 22312 12000 22432 6 wbm_a_adr_o[22]
port 19 nsew signal tristate
rlabel metal3 s 11200 23128 12000 23248 6 wbm_a_adr_o[23]
port 20 nsew signal tristate
rlabel metal3 s 11200 23808 12000 23928 6 wbm_a_adr_o[24]
port 21 nsew signal tristate
rlabel metal3 s 11200 24624 12000 24744 6 wbm_a_adr_o[25]
port 22 nsew signal tristate
rlabel metal3 s 11200 25304 12000 25424 6 wbm_a_adr_o[26]
port 23 nsew signal tristate
rlabel metal3 s 11200 26120 12000 26240 6 wbm_a_adr_o[27]
port 24 nsew signal tristate
rlabel metal3 s 11200 26936 12000 27056 6 wbm_a_adr_o[28]
port 25 nsew signal tristate
rlabel metal3 s 11200 27616 12000 27736 6 wbm_a_adr_o[29]
port 26 nsew signal tristate
rlabel metal3 s 11200 7080 12000 7200 6 wbm_a_adr_o[2]
port 27 nsew signal tristate
rlabel metal3 s 11200 28432 12000 28552 6 wbm_a_adr_o[30]
port 28 nsew signal tristate
rlabel metal3 s 11200 29112 12000 29232 6 wbm_a_adr_o[31]
port 29 nsew signal tristate
rlabel metal3 s 11200 7896 12000 8016 6 wbm_a_adr_o[3]
port 30 nsew signal tristate
rlabel metal3 s 11200 8576 12000 8696 6 wbm_a_adr_o[4]
port 31 nsew signal tristate
rlabel metal3 s 11200 9392 12000 9512 6 wbm_a_adr_o[5]
port 32 nsew signal tristate
rlabel metal3 s 11200 10072 12000 10192 6 wbm_a_adr_o[6]
port 33 nsew signal tristate
rlabel metal3 s 11200 10888 12000 11008 6 wbm_a_adr_o[7]
port 34 nsew signal tristate
rlabel metal3 s 11200 11704 12000 11824 6 wbm_a_adr_o[8]
port 35 nsew signal tristate
rlabel metal3 s 11200 12384 12000 12504 6 wbm_a_adr_o[9]
port 36 nsew signal tristate
rlabel metal3 s 11200 960 12000 1080 6 wbm_a_cyc_o
port 37 nsew signal tristate
rlabel metal3 s 11200 54272 12000 54392 6 wbm_a_dat_i[0]
port 38 nsew signal input
rlabel metal3 s 11200 61888 12000 62008 6 wbm_a_dat_i[10]
port 39 nsew signal input
rlabel metal3 s 11200 62704 12000 62824 6 wbm_a_dat_i[11]
port 40 nsew signal input
rlabel metal3 s 11200 63384 12000 63504 6 wbm_a_dat_i[12]
port 41 nsew signal input
rlabel metal3 s 11200 64200 12000 64320 6 wbm_a_dat_i[13]
port 42 nsew signal input
rlabel metal3 s 11200 65016 12000 65136 6 wbm_a_dat_i[14]
port 43 nsew signal input
rlabel metal3 s 11200 65696 12000 65816 6 wbm_a_dat_i[15]
port 44 nsew signal input
rlabel metal3 s 11200 66512 12000 66632 6 wbm_a_dat_i[16]
port 45 nsew signal input
rlabel metal3 s 11200 67192 12000 67312 6 wbm_a_dat_i[17]
port 46 nsew signal input
rlabel metal3 s 11200 68008 12000 68128 6 wbm_a_dat_i[18]
port 47 nsew signal input
rlabel metal3 s 11200 68824 12000 68944 6 wbm_a_dat_i[19]
port 48 nsew signal input
rlabel metal3 s 11200 55088 12000 55208 6 wbm_a_dat_i[1]
port 49 nsew signal input
rlabel metal3 s 11200 69504 12000 69624 6 wbm_a_dat_i[20]
port 50 nsew signal input
rlabel metal3 s 11200 70320 12000 70440 6 wbm_a_dat_i[21]
port 51 nsew signal input
rlabel metal3 s 11200 71000 12000 71120 6 wbm_a_dat_i[22]
port 52 nsew signal input
rlabel metal3 s 11200 71816 12000 71936 6 wbm_a_dat_i[23]
port 53 nsew signal input
rlabel metal3 s 11200 72632 12000 72752 6 wbm_a_dat_i[24]
port 54 nsew signal input
rlabel metal3 s 11200 73312 12000 73432 6 wbm_a_dat_i[25]
port 55 nsew signal input
rlabel metal3 s 11200 74128 12000 74248 6 wbm_a_dat_i[26]
port 56 nsew signal input
rlabel metal3 s 11200 74808 12000 74928 6 wbm_a_dat_i[27]
port 57 nsew signal input
rlabel metal3 s 11200 75624 12000 75744 6 wbm_a_dat_i[28]
port 58 nsew signal input
rlabel metal3 s 11200 76440 12000 76560 6 wbm_a_dat_i[29]
port 59 nsew signal input
rlabel metal3 s 11200 55768 12000 55888 6 wbm_a_dat_i[2]
port 60 nsew signal input
rlabel metal3 s 11200 77120 12000 77240 6 wbm_a_dat_i[30]
port 61 nsew signal input
rlabel metal3 s 11200 77936 12000 78056 6 wbm_a_dat_i[31]
port 62 nsew signal input
rlabel metal3 s 11200 56584 12000 56704 6 wbm_a_dat_i[3]
port 63 nsew signal input
rlabel metal3 s 11200 57400 12000 57520 6 wbm_a_dat_i[4]
port 64 nsew signal input
rlabel metal3 s 11200 58080 12000 58200 6 wbm_a_dat_i[5]
port 65 nsew signal input
rlabel metal3 s 11200 58896 12000 59016 6 wbm_a_dat_i[6]
port 66 nsew signal input
rlabel metal3 s 11200 59576 12000 59696 6 wbm_a_dat_i[7]
port 67 nsew signal input
rlabel metal3 s 11200 60392 12000 60512 6 wbm_a_dat_i[8]
port 68 nsew signal input
rlabel metal3 s 11200 61208 12000 61328 6 wbm_a_dat_i[9]
port 69 nsew signal input
rlabel metal3 s 11200 29928 12000 30048 6 wbm_a_dat_o[0]
port 70 nsew signal tristate
rlabel metal3 s 11200 37544 12000 37664 6 wbm_a_dat_o[10]
port 71 nsew signal tristate
rlabel metal3 s 11200 38360 12000 38480 6 wbm_a_dat_o[11]
port 72 nsew signal tristate
rlabel metal3 s 11200 39040 12000 39160 6 wbm_a_dat_o[12]
port 73 nsew signal tristate
rlabel metal3 s 11200 39856 12000 39976 6 wbm_a_dat_o[13]
port 74 nsew signal tristate
rlabel metal3 s 11200 40536 12000 40656 6 wbm_a_dat_o[14]
port 75 nsew signal tristate
rlabel metal3 s 11200 41352 12000 41472 6 wbm_a_dat_o[15]
port 76 nsew signal tristate
rlabel metal3 s 11200 42168 12000 42288 6 wbm_a_dat_o[16]
port 77 nsew signal tristate
rlabel metal3 s 11200 42848 12000 42968 6 wbm_a_dat_o[17]
port 78 nsew signal tristate
rlabel metal3 s 11200 43664 12000 43784 6 wbm_a_dat_o[18]
port 79 nsew signal tristate
rlabel metal3 s 11200 44344 12000 44464 6 wbm_a_dat_o[19]
port 80 nsew signal tristate
rlabel metal3 s 11200 30744 12000 30864 6 wbm_a_dat_o[1]
port 81 nsew signal tristate
rlabel metal3 s 11200 45160 12000 45280 6 wbm_a_dat_o[20]
port 82 nsew signal tristate
rlabel metal3 s 11200 45976 12000 46096 6 wbm_a_dat_o[21]
port 83 nsew signal tristate
rlabel metal3 s 11200 46656 12000 46776 6 wbm_a_dat_o[22]
port 84 nsew signal tristate
rlabel metal3 s 11200 47472 12000 47592 6 wbm_a_dat_o[23]
port 85 nsew signal tristate
rlabel metal3 s 11200 48152 12000 48272 6 wbm_a_dat_o[24]
port 86 nsew signal tristate
rlabel metal3 s 11200 48968 12000 49088 6 wbm_a_dat_o[25]
port 87 nsew signal tristate
rlabel metal3 s 11200 49784 12000 49904 6 wbm_a_dat_o[26]
port 88 nsew signal tristate
rlabel metal3 s 11200 50464 12000 50584 6 wbm_a_dat_o[27]
port 89 nsew signal tristate
rlabel metal3 s 11200 51280 12000 51400 6 wbm_a_dat_o[28]
port 90 nsew signal tristate
rlabel metal3 s 11200 51960 12000 52080 6 wbm_a_dat_o[29]
port 91 nsew signal tristate
rlabel metal3 s 11200 31424 12000 31544 6 wbm_a_dat_o[2]
port 92 nsew signal tristate
rlabel metal3 s 11200 52776 12000 52896 6 wbm_a_dat_o[30]
port 93 nsew signal tristate
rlabel metal3 s 11200 53592 12000 53712 6 wbm_a_dat_o[31]
port 94 nsew signal tristate
rlabel metal3 s 11200 32240 12000 32360 6 wbm_a_dat_o[3]
port 95 nsew signal tristate
rlabel metal3 s 11200 32920 12000 33040 6 wbm_a_dat_o[4]
port 96 nsew signal tristate
rlabel metal3 s 11200 33736 12000 33856 6 wbm_a_dat_o[5]
port 97 nsew signal tristate
rlabel metal3 s 11200 34552 12000 34672 6 wbm_a_dat_o[6]
port 98 nsew signal tristate
rlabel metal3 s 11200 35232 12000 35352 6 wbm_a_dat_o[7]
port 99 nsew signal tristate
rlabel metal3 s 11200 36048 12000 36168 6 wbm_a_dat_o[8]
port 100 nsew signal tristate
rlabel metal3 s 11200 36728 12000 36848 6 wbm_a_dat_o[9]
port 101 nsew signal tristate
rlabel metal3 s 11200 2456 12000 2576 6 wbm_a_sel_o[0]
port 102 nsew signal tristate
rlabel metal3 s 11200 3272 12000 3392 6 wbm_a_sel_o[1]
port 103 nsew signal tristate
rlabel metal3 s 11200 4088 12000 4208 6 wbm_a_sel_o[2]
port 104 nsew signal tristate
rlabel metal3 s 11200 4768 12000 4888 6 wbm_a_sel_o[3]
port 105 nsew signal tristate
rlabel metal3 s 11200 280 12000 400 6 wbm_a_stb_o
port 106 nsew signal tristate
rlabel metal3 s 11200 1776 12000 1896 6 wbm_a_we_o
port 107 nsew signal tristate
rlabel metal3 s 0 79568 800 79688 6 wbm_b_ack_i
port 108 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 wbm_b_adr_o[0]
port 109 nsew signal tristate
rlabel metal3 s 0 48288 800 48408 6 wbm_b_adr_o[1]
port 110 nsew signal tristate
rlabel metal3 s 0 48696 800 48816 6 wbm_b_adr_o[2]
port 111 nsew signal tristate
rlabel metal3 s 0 49104 800 49224 6 wbm_b_adr_o[3]
port 112 nsew signal tristate
rlabel metal3 s 0 49512 800 49632 6 wbm_b_adr_o[4]
port 113 nsew signal tristate
rlabel metal3 s 0 49920 800 50040 6 wbm_b_adr_o[5]
port 114 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 wbm_b_adr_o[6]
port 115 nsew signal tristate
rlabel metal3 s 0 50872 800 50992 6 wbm_b_adr_o[7]
port 116 nsew signal tristate
rlabel metal3 s 0 51280 800 51400 6 wbm_b_adr_o[8]
port 117 nsew signal tristate
rlabel metal3 s 0 51688 800 51808 6 wbm_b_adr_o[9]
port 118 nsew signal tristate
rlabel metal3 s 0 45160 800 45280 6 wbm_b_cyc_o
port 119 nsew signal tristate
rlabel metal3 s 0 65832 800 65952 6 wbm_b_dat_i[0]
port 120 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbm_b_dat_i[10]
port 121 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 wbm_b_dat_i[11]
port 122 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 wbm_b_dat_i[12]
port 123 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 wbm_b_dat_i[13]
port 124 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 wbm_b_dat_i[14]
port 125 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbm_b_dat_i[15]
port 126 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 wbm_b_dat_i[16]
port 127 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 wbm_b_dat_i[17]
port 128 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 wbm_b_dat_i[18]
port 129 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 wbm_b_dat_i[19]
port 130 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 wbm_b_dat_i[1]
port 131 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 wbm_b_dat_i[20]
port 132 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 wbm_b_dat_i[21]
port 133 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 wbm_b_dat_i[22]
port 134 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 wbm_b_dat_i[23]
port 135 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 wbm_b_dat_i[24]
port 136 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 wbm_b_dat_i[25]
port 137 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 wbm_b_dat_i[26]
port 138 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 wbm_b_dat_i[27]
port 139 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 wbm_b_dat_i[28]
port 140 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 wbm_b_dat_i[29]
port 141 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 wbm_b_dat_i[2]
port 142 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 wbm_b_dat_i[30]
port 143 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 wbm_b_dat_i[31]
port 144 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 wbm_b_dat_i[3]
port 145 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 wbm_b_dat_i[4]
port 146 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 wbm_b_dat_i[5]
port 147 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 wbm_b_dat_i[6]
port 148 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 wbm_b_dat_i[7]
port 149 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wbm_b_dat_i[8]
port 150 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 wbm_b_dat_i[9]
port 151 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 wbm_b_dat_o[0]
port 152 nsew signal tristate
rlabel metal3 s 0 56448 800 56568 6 wbm_b_dat_o[10]
port 153 nsew signal tristate
rlabel metal3 s 0 56856 800 56976 6 wbm_b_dat_o[11]
port 154 nsew signal tristate
rlabel metal3 s 0 57264 800 57384 6 wbm_b_dat_o[12]
port 155 nsew signal tristate
rlabel metal3 s 0 57672 800 57792 6 wbm_b_dat_o[13]
port 156 nsew signal tristate
rlabel metal3 s 0 58080 800 58200 6 wbm_b_dat_o[14]
port 157 nsew signal tristate
rlabel metal3 s 0 58488 800 58608 6 wbm_b_dat_o[15]
port 158 nsew signal tristate
rlabel metal3 s 0 59032 800 59152 6 wbm_b_dat_o[16]
port 159 nsew signal tristate
rlabel metal3 s 0 59440 800 59560 6 wbm_b_dat_o[17]
port 160 nsew signal tristate
rlabel metal3 s 0 59848 800 59968 6 wbm_b_dat_o[18]
port 161 nsew signal tristate
rlabel metal3 s 0 60256 800 60376 6 wbm_b_dat_o[19]
port 162 nsew signal tristate
rlabel metal3 s 0 52504 800 52624 6 wbm_b_dat_o[1]
port 163 nsew signal tristate
rlabel metal3 s 0 60664 800 60784 6 wbm_b_dat_o[20]
port 164 nsew signal tristate
rlabel metal3 s 0 61072 800 61192 6 wbm_b_dat_o[21]
port 165 nsew signal tristate
rlabel metal3 s 0 61616 800 61736 6 wbm_b_dat_o[22]
port 166 nsew signal tristate
rlabel metal3 s 0 62024 800 62144 6 wbm_b_dat_o[23]
port 167 nsew signal tristate
rlabel metal3 s 0 62432 800 62552 6 wbm_b_dat_o[24]
port 168 nsew signal tristate
rlabel metal3 s 0 62840 800 62960 6 wbm_b_dat_o[25]
port 169 nsew signal tristate
rlabel metal3 s 0 63248 800 63368 6 wbm_b_dat_o[26]
port 170 nsew signal tristate
rlabel metal3 s 0 63656 800 63776 6 wbm_b_dat_o[27]
port 171 nsew signal tristate
rlabel metal3 s 0 64200 800 64320 6 wbm_b_dat_o[28]
port 172 nsew signal tristate
rlabel metal3 s 0 64608 800 64728 6 wbm_b_dat_o[29]
port 173 nsew signal tristate
rlabel metal3 s 0 52912 800 53032 6 wbm_b_dat_o[2]
port 174 nsew signal tristate
rlabel metal3 s 0 65016 800 65136 6 wbm_b_dat_o[30]
port 175 nsew signal tristate
rlabel metal3 s 0 65424 800 65544 6 wbm_b_dat_o[31]
port 176 nsew signal tristate
rlabel metal3 s 0 53456 800 53576 6 wbm_b_dat_o[3]
port 177 nsew signal tristate
rlabel metal3 s 0 53864 800 53984 6 wbm_b_dat_o[4]
port 178 nsew signal tristate
rlabel metal3 s 0 54272 800 54392 6 wbm_b_dat_o[5]
port 179 nsew signal tristate
rlabel metal3 s 0 54680 800 54800 6 wbm_b_dat_o[6]
port 180 nsew signal tristate
rlabel metal3 s 0 55088 800 55208 6 wbm_b_dat_o[7]
port 181 nsew signal tristate
rlabel metal3 s 0 55496 800 55616 6 wbm_b_dat_o[8]
port 182 nsew signal tristate
rlabel metal3 s 0 55904 800 56024 6 wbm_b_dat_o[9]
port 183 nsew signal tristate
rlabel metal3 s 0 46112 800 46232 6 wbm_b_sel_o[0]
port 184 nsew signal tristate
rlabel metal3 s 0 46520 800 46640 6 wbm_b_sel_o[1]
port 185 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 wbm_b_sel_o[2]
port 186 nsew signal tristate
rlabel metal3 s 0 47336 800 47456 6 wbm_b_sel_o[3]
port 187 nsew signal tristate
rlabel metal3 s 0 44752 800 44872 6 wbm_b_stb_o
port 188 nsew signal tristate
rlabel metal3 s 0 45704 800 45824 6 wbm_b_we_o
port 189 nsew signal tristate
rlabel metal3 s 0 44344 800 44464 6 wbs_ack_o
port 190 nsew signal tristate
rlabel metal3 s 0 3136 800 3256 6 wbs_adr_i[0]
port 191 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 wbs_adr_i[10]
port 192 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 wbs_adr_i[11]
port 193 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 wbs_adr_i[12]
port 194 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 wbs_adr_i[13]
port 195 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 wbs_adr_i[14]
port 196 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wbs_adr_i[15]
port 197 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 wbs_adr_i[16]
port 198 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 wbs_adr_i[17]
port 199 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_adr_i[18]
port 200 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 wbs_adr_i[19]
port 201 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 wbs_adr_i[1]
port 202 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 wbs_adr_i[20]
port 203 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 wbs_adr_i[21]
port 204 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 wbs_adr_i[22]
port 205 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_adr_i[23]
port 206 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 wbs_adr_i[24]
port 207 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 wbs_adr_i[25]
port 208 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 wbs_adr_i[26]
port 209 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 wbs_adr_i[27]
port 210 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 wbs_adr_i[28]
port 211 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 wbs_adr_i[29]
port 212 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 wbs_adr_i[2]
port 213 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 wbs_adr_i[30]
port 214 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 wbs_adr_i[31]
port 215 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 wbs_adr_i[3]
port 216 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wbs_adr_i[4]
port 217 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 wbs_adr_i[5]
port 218 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 wbs_adr_i[6]
port 219 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wbs_adr_i[7]
port 220 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 wbs_adr_i[8]
port 221 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 wbs_adr_i[9]
port 222 nsew signal input
rlabel metal3 s 0 552 800 672 6 wbs_cyc_i
port 223 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 wbs_dat_i[0]
port 224 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_i[10]
port 225 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 wbs_dat_i[11]
port 226 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 wbs_dat_i[12]
port 227 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wbs_dat_i[13]
port 228 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 wbs_dat_i[14]
port 229 nsew signal input
rlabel metal3 s 0 23264 800 23384 6 wbs_dat_i[15]
port 230 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 wbs_dat_i[16]
port 231 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 wbs_dat_i[17]
port 232 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 wbs_dat_i[18]
port 233 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 wbs_dat_i[19]
port 234 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 wbs_dat_i[1]
port 235 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 wbs_dat_i[20]
port 236 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_dat_i[21]
port 237 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 wbs_dat_i[22]
port 238 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 wbs_dat_i[23]
port 239 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wbs_dat_i[24]
port 240 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 wbs_dat_i[25]
port 241 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 wbs_dat_i[26]
port 242 nsew signal input
rlabel metal3 s 0 28432 800 28552 6 wbs_dat_i[27]
port 243 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 wbs_dat_i[28]
port 244 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_i[29]
port 245 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 wbs_dat_i[2]
port 246 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 wbs_dat_i[30]
port 247 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 wbs_dat_i[31]
port 248 nsew signal input
rlabel metal3 s 0 18096 800 18216 6 wbs_dat_i[3]
port 249 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 wbs_dat_i[4]
port 250 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wbs_dat_i[5]
port 251 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 wbs_dat_i[6]
port 252 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 wbs_dat_i[7]
port 253 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wbs_dat_i[8]
port 254 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 wbs_dat_i[9]
port 255 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 wbs_dat_o[0]
port 256 nsew signal tristate
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_o[10]
port 257 nsew signal tristate
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_o[11]
port 258 nsew signal tristate
rlabel metal3 s 0 35776 800 35896 6 wbs_dat_o[12]
port 259 nsew signal tristate
rlabel metal3 s 0 36184 800 36304 6 wbs_dat_o[13]
port 260 nsew signal tristate
rlabel metal3 s 0 36592 800 36712 6 wbs_dat_o[14]
port 261 nsew signal tristate
rlabel metal3 s 0 37000 800 37120 6 wbs_dat_o[15]
port 262 nsew signal tristate
rlabel metal3 s 0 37544 800 37664 6 wbs_dat_o[16]
port 263 nsew signal tristate
rlabel metal3 s 0 37952 800 38072 6 wbs_dat_o[17]
port 264 nsew signal tristate
rlabel metal3 s 0 38360 800 38480 6 wbs_dat_o[18]
port 265 nsew signal tristate
rlabel metal3 s 0 38768 800 38888 6 wbs_dat_o[19]
port 266 nsew signal tristate
rlabel metal3 s 0 31016 800 31136 6 wbs_dat_o[1]
port 267 nsew signal tristate
rlabel metal3 s 0 39176 800 39296 6 wbs_dat_o[20]
port 268 nsew signal tristate
rlabel metal3 s 0 39584 800 39704 6 wbs_dat_o[21]
port 269 nsew signal tristate
rlabel metal3 s 0 40128 800 40248 6 wbs_dat_o[22]
port 270 nsew signal tristate
rlabel metal3 s 0 40536 800 40656 6 wbs_dat_o[23]
port 271 nsew signal tristate
rlabel metal3 s 0 40944 800 41064 6 wbs_dat_o[24]
port 272 nsew signal tristate
rlabel metal3 s 0 41352 800 41472 6 wbs_dat_o[25]
port 273 nsew signal tristate
rlabel metal3 s 0 41760 800 41880 6 wbs_dat_o[26]
port 274 nsew signal tristate
rlabel metal3 s 0 42168 800 42288 6 wbs_dat_o[27]
port 275 nsew signal tristate
rlabel metal3 s 0 42576 800 42696 6 wbs_dat_o[28]
port 276 nsew signal tristate
rlabel metal3 s 0 43120 800 43240 6 wbs_dat_o[29]
port 277 nsew signal tristate
rlabel metal3 s 0 31424 800 31544 6 wbs_dat_o[2]
port 278 nsew signal tristate
rlabel metal3 s 0 43528 800 43648 6 wbs_dat_o[30]
port 279 nsew signal tristate
rlabel metal3 s 0 43936 800 44056 6 wbs_dat_o[31]
port 280 nsew signal tristate
rlabel metal3 s 0 31832 800 31952 6 wbs_dat_o[3]
port 281 nsew signal tristate
rlabel metal3 s 0 32376 800 32496 6 wbs_dat_o[4]
port 282 nsew signal tristate
rlabel metal3 s 0 32784 800 32904 6 wbs_dat_o[5]
port 283 nsew signal tristate
rlabel metal3 s 0 33192 800 33312 6 wbs_dat_o[6]
port 284 nsew signal tristate
rlabel metal3 s 0 33600 800 33720 6 wbs_dat_o[7]
port 285 nsew signal tristate
rlabel metal3 s 0 34008 800 34128 6 wbs_dat_o[8]
port 286 nsew signal tristate
rlabel metal3 s 0 34416 800 34536 6 wbs_dat_o[9]
port 287 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 wbs_sel_i[0]
port 288 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 wbs_sel_i[1]
port 289 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 wbs_sel_i[2]
port 290 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 wbs_sel_i[3]
port 291 nsew signal input
rlabel metal3 s 0 144 800 264 6 wbs_stb_i
port 292 nsew signal input
rlabel metal3 s 0 960 800 1080 6 wbs_we_i
port 293 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 12000 80000
<< end >>
